/*
 * Copyright (c) 2025 ROOTS Education Co.
 * based on the VGA examples by Uri Shaked
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

parameter LOGO_SIZE = 256;  // Size of the logo in pixels
parameter DISPLAY_WIDTH = 640;  // VGA display width
parameter DISPLAY_HEIGHT = 480;  // VGA display height

`define COLOR_WHITE 3'd7

module tt_um_arud4172_ROOTS_vga (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;

  // Configuration
  wire cfg_tile = ui_in[0];
  wire cfg_color = ui_in[1];

  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  reg [9:0] prev_y;

  hvsync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );

  reg [9:0] logo_left;
  reg [9:0] logo_top;
  reg dir_x;
  reg dir_y;

  wire pixel_value;
  reg [2:0] color_index;
  wire [5:0] color;

  wire [9:0] x = pix_x - logo_left;
  wire [9:0] y = pix_y - logo_top;
  wire logo_pixels = cfg_tile || (x < LOGO_SIZE && y < LOGO_SIZE);

  bitmap_rom rom1 (
      .x(x[7:0]),
      .y(y[7:0]),
      .pixel(pixel_value)
  );

  palette palette_inst (
      .color_index(cfg_color ? color_index : `COLOR_WHITE),
      .rrggbb(color)
  );

  // RGB output logic

  reg [7:0] frame_counter;

  // Mirror pixel positions to create kaleidoscope symmetry
  // Original animation (fast)
  wire [9:0] mx = (pix_x + frame_counter) ^ (pix_y >> 1);
  wire [9:0] my = (pix_y + frame_counter) ^ (pix_x >> 1);

  // Generate pattern
  wire kaleido_bit = mx[5] ^ my[5];  // 32-pixel symmetric pattern

  // Create some color shifting
  wire [1:0] kaleido_r = mx[7:6];
  wire [1:0] kaleido_g = my[7:6];
  wire [1:0] kaleido_b = {mx[6] ^ my[6], mx[5] ^ my[5]};

  always @(posedge clk) begin
    if (~rst_n) begin
      R <= 0;
      G <= 0;
      B <= 0;
    end else begin
      R <= 0;
      G <= 0;
      B <= 0;

      if (video_active) begin
        if (logo_pixels && pixel_value) begin
          // Foreground logo
          R <= color[5:4];
          G <= color[3:2];
          B <= color[1:0];
        end else begin
          // Kaleidoscope background
          R <= kaleido_bit ? kaleido_r : ~kaleido_r;
          G <= kaleido_bit ? kaleido_g : ~kaleido_g;
          B <= kaleido_bit ? kaleido_b : ~kaleido_b;
        end
      end
    end
  end


  // Bouncing logic
  always @(posedge clk) begin
    if (~rst_n) begin
      logo_left <= (DISPLAY_WIDTH - LOGO_SIZE) / 2;
      logo_top  <= (DISPLAY_HEIGHT - LOGO_SIZE) / 2;
      dir_y <= 0;
      dir_x <= 1;
      color_index <= 0;
    end else begin
      prev_y <= pix_y;
      if (pix_y == 0 && prev_y != pix_y) begin
        logo_left <= logo_left + (dir_x ? 1 : -1);
        logo_top  <= logo_top + (dir_y ? 1 : -1);
        frame_counter <= frame_counter + 1;
        if (logo_left - 1 == 0 && !dir_x) begin
          dir_x <= 1;
          color_index <= color_index + 1;
        end
        if (logo_left + 1 >= DISPLAY_WIDTH - LOGO_SIZE && dir_x) begin
          dir_x <= 0;
          color_index <= color_index + 1;
        end
        if (logo_top - 1 == 0 && !dir_y) begin
          dir_y <= 1;
          color_index <= color_index + 1;
        end
        if (logo_top + 1 == DISPLAY_HEIGHT - LOGO_SIZE && dir_y) begin
          dir_y <= 0;
          color_index <= color_index + 1;
        end
      end
    end
  end

endmodule

`default_nettype none

/*
Video sync generator, used to drive a VGA monitor.
Timing from: https://en.wikipedia.org/wiki/Video_Graphics_Array
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
*/

module vga_sync_generator (
    clk,
    reset,
    hsync,
    vsync,
    display_on,
    hpos,
    vpos
);

  input clk;
  input reset;
  output reg hsync, vsync;
  output display_on;
  output reg [9:0] hpos;
  output reg [9:0] vpos;

  // declarations for TV-simulator sync parameters
  // horizontal constants
  parameter H_DISPLAY = 640;  // horizontal display width
  parameter H_BACK = 48;  // horizontal left border (back porch)
  parameter H_FRONT = 16;  // horizontal right border (front porch)
  parameter H_SYNC = 96;  // horizontal sync width
  // vertical constants
  parameter V_DISPLAY = 480;  // vertical display height
  parameter V_TOP = 33;  // vertical top border
  parameter V_BOTTOM = 10;  // vertical bottom border
  parameter V_SYNC = 2;  // vertical sync # lines
  // derived constants
  parameter H_SYNC_START = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START = V_DISPLAY + V_BOTTOM;
  parameter V_SYNC_END = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
  parameter V_MAX = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

  wire hmaxxed = (hpos == H_MAX) || reset;  // set when hpos is maximum
  wire vmaxxed = (vpos == V_MAX) || reset;  // set when vpos is maximum

  // horizontal position counter
  always @(posedge clk) begin
    hsync <= (hpos >= H_SYNC_START && hpos <= H_SYNC_END);
    if (hmaxxed) hpos <= 0;
    else hpos <= hpos + 1;
  end

  // vertical position counter
  always @(posedge clk) begin
    vsync <= (vpos >= V_SYNC_START && vpos <= V_SYNC_END);
    if (hmaxxed)
      if (vmaxxed) vpos <= 0;
      else vpos <= vpos + 1;
  end

  // display_on is set when beam is in "safe" visible frame
  assign display_on = (hpos < H_DISPLAY) && (vpos < V_DISPLAY);

endmodule

// --------------------------------------------------------

module palette (
    input  wire [2:0] color_index,
    output wire [5:0] rrggbb
);

  reg [5:0] palette[7:0];

  initial begin
    palette[0] = 6'b001011;  // cyan
    palette[1] = 6'b110110;  // pink
    palette[2] = 6'b101101;  // green
    palette[3] = 6'b111000;  // orange
    palette[4] = 6'b110011;  // purple
    palette[5] = 6'b011111;  // yellow 
    palette[6] = 6'b110001;  // red
    palette[7] = 6'b111111;  // white
  end

  assign rrggbb = palette[color_index];

endmodule

// --------------------------------------------------------

module bitmap_rom (
    input wire [7:0] x,
    input wire [7:0] y,
    output wire pixel
);
  reg [7:0] mem[8191:0];  // 256 rows × 32 bytes = 8192 bytes

  wire [12:0] addr = (y << 5) + (x >> 3);  // y * 32 + x / 8
  assign pixel = mem[addr][7 - x[2:0]];

  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'h00;
    mem[164] = 8'h00;
    mem[165] = 8'h00;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'h00;
    mem[171] = 8'h00;
    mem[172] = 8'h00;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'h00;
    mem[180] = 8'h00;
    mem[181] = 8'h00;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'h00;
    mem[187] = 8'h00;
    mem[188] = 8'h00;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'h00;
    mem[195] = 8'h00;
    mem[196] = 8'h00;
    mem[197] = 8'h00;
    mem[198] = 8'h00;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'h00;
    mem[202] = 8'h00;
    mem[203] = 8'h00;
    mem[204] = 8'h00;
    mem[205] = 8'h00;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'h00;
    mem[211] = 8'h00;
    mem[212] = 8'h00;
    mem[213] = 8'h00;
    mem[214] = 8'h00;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'h00;
    mem[219] = 8'h00;
    mem[220] = 8'h00;
    mem[221] = 8'h00;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h00;
    mem[227] = 8'h00;
    mem[228] = 8'h00;
    mem[229] = 8'h00;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h00;
    mem[235] = 8'h00;
    mem[236] = 8'h00;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h00;
    mem[243] = 8'h00;
    mem[244] = 8'h00;
    mem[245] = 8'h00;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'h00;
    mem[251] = 8'h00;
    mem[252] = 8'h00;
    mem[253] = 8'h00;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'h00;
    mem[259] = 8'h00;
    mem[260] = 8'h00;
    mem[261] = 8'h00;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'h00;
    mem[267] = 8'h00;
    mem[268] = 8'h00;
    mem[269] = 8'h00;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'h00;
    mem[275] = 8'h00;
    mem[276] = 8'h00;
    mem[277] = 8'h00;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h00;
    mem[283] = 8'h00;
    mem[284] = 8'h00;
    mem[285] = 8'h00;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'h00;
    mem[291] = 8'h00;
    mem[292] = 8'h00;
    mem[293] = 8'h00;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'h00;
    mem[300] = 8'h00;
    mem[301] = 8'h00;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'h00;
    mem[307] = 8'h00;
    mem[308] = 8'h00;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'h00;
    mem[316] = 8'h00;
    mem[317] = 8'h00;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'h00;
    mem[323] = 8'h00;
    mem[324] = 8'h00;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'h00;
    mem[332] = 8'h00;
    mem[333] = 8'h00;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'h00;
    mem[339] = 8'h00;
    mem[340] = 8'h00;
    mem[341] = 8'h00;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'h00;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'h00;
    mem[355] = 8'h00;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'hf0;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'hfe;
    mem[432] = 8'h03;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h80;
    mem[463] = 8'hff;
    mem[464] = 8'h1f;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'he0;
    mem[495] = 8'hff;
    mem[496] = 8'h7f;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
    mem[512] = 8'h00;
    mem[513] = 8'h00;
    mem[514] = 8'h00;
    mem[515] = 8'h00;
    mem[516] = 8'h00;
    mem[517] = 8'h00;
    mem[518] = 8'h00;
    mem[519] = 8'h00;
    mem[520] = 8'h00;
    mem[521] = 8'h00;
    mem[522] = 8'h00;
    mem[523] = 8'h00;
    mem[524] = 8'h00;
    mem[525] = 8'h00;
    mem[526] = 8'hf8;
    mem[527] = 8'hff;
    mem[528] = 8'hff;
    mem[529] = 8'h01;
    mem[530] = 8'h00;
    mem[531] = 8'h00;
    mem[532] = 8'h00;
    mem[533] = 8'h00;
    mem[534] = 8'h00;
    mem[535] = 8'h00;
    mem[536] = 8'h00;
    mem[537] = 8'h00;
    mem[538] = 8'h00;
    mem[539] = 8'h00;
    mem[540] = 8'h00;
    mem[541] = 8'h00;
    mem[542] = 8'h00;
    mem[543] = 8'h00;
    mem[544] = 8'h00;
    mem[545] = 8'h00;
    mem[546] = 8'h00;
    mem[547] = 8'h00;
    mem[548] = 8'h00;
    mem[549] = 8'h00;
    mem[550] = 8'h00;
    mem[551] = 8'h00;
    mem[552] = 8'h00;
    mem[553] = 8'h00;
    mem[554] = 8'h00;
    mem[555] = 8'h00;
    mem[556] = 8'h00;
    mem[557] = 8'h00;
    mem[558] = 8'hfe;
    mem[559] = 8'hff;
    mem[560] = 8'hff;
    mem[561] = 8'h07;
    mem[562] = 8'h00;
    mem[563] = 8'h00;
    mem[564] = 8'h00;
    mem[565] = 8'h00;
    mem[566] = 8'h00;
    mem[567] = 8'h00;
    mem[568] = 8'h00;
    mem[569] = 8'h00;
    mem[570] = 8'h00;
    mem[571] = 8'h00;
    mem[572] = 8'h00;
    mem[573] = 8'h00;
    mem[574] = 8'h00;
    mem[575] = 8'h00;
    mem[576] = 8'h00;
    mem[577] = 8'h00;
    mem[578] = 8'h00;
    mem[579] = 8'h00;
    mem[580] = 8'h00;
    mem[581] = 8'h00;
    mem[582] = 8'h00;
    mem[583] = 8'h00;
    mem[584] = 8'h00;
    mem[585] = 8'h00;
    mem[586] = 8'h00;
    mem[587] = 8'h00;
    mem[588] = 8'h00;
    mem[589] = 8'h80;
    mem[590] = 8'hff;
    mem[591] = 8'hff;
    mem[592] = 8'hff;
    mem[593] = 8'h1f;
    mem[594] = 8'h00;
    mem[595] = 8'h00;
    mem[596] = 8'h00;
    mem[597] = 8'h00;
    mem[598] = 8'h00;
    mem[599] = 8'h00;
    mem[600] = 8'h00;
    mem[601] = 8'h00;
    mem[602] = 8'h00;
    mem[603] = 8'h00;
    mem[604] = 8'h00;
    mem[605] = 8'h00;
    mem[606] = 8'h00;
    mem[607] = 8'h00;
    mem[608] = 8'h00;
    mem[609] = 8'h00;
    mem[610] = 8'h00;
    mem[611] = 8'h00;
    mem[612] = 8'h00;
    mem[613] = 8'h00;
    mem[614] = 8'h00;
    mem[615] = 8'h00;
    mem[616] = 8'h00;
    mem[617] = 8'h00;
    mem[618] = 8'h00;
    mem[619] = 8'h00;
    mem[620] = 8'h00;
    mem[621] = 8'he0;
    mem[622] = 8'hff;
    mem[623] = 8'hff;
    mem[624] = 8'hff;
    mem[625] = 8'h7f;
    mem[626] = 8'h00;
    mem[627] = 8'h00;
    mem[628] = 8'h00;
    mem[629] = 8'h00;
    mem[630] = 8'h00;
    mem[631] = 8'h00;
    mem[632] = 8'h00;
    mem[633] = 8'h00;
    mem[634] = 8'h00;
    mem[635] = 8'h00;
    mem[636] = 8'h00;
    mem[637] = 8'h00;
    mem[638] = 8'h00;
    mem[639] = 8'h00;
    mem[640] = 8'h00;
    mem[641] = 8'h00;
    mem[642] = 8'h00;
    mem[643] = 8'h00;
    mem[644] = 8'h00;
    mem[645] = 8'h00;
    mem[646] = 8'h00;
    mem[647] = 8'h00;
    mem[648] = 8'h00;
    mem[649] = 8'h00;
    mem[650] = 8'h00;
    mem[651] = 8'h00;
    mem[652] = 8'h00;
    mem[653] = 8'hf8;
    mem[654] = 8'hff;
    mem[655] = 8'h0f;
    mem[656] = 8'hff;
    mem[657] = 8'hff;
    mem[658] = 8'h01;
    mem[659] = 8'h00;
    mem[660] = 8'h00;
    mem[661] = 8'h00;
    mem[662] = 8'h00;
    mem[663] = 8'h00;
    mem[664] = 8'h00;
    mem[665] = 8'h00;
    mem[666] = 8'h00;
    mem[667] = 8'h00;
    mem[668] = 8'h00;
    mem[669] = 8'h00;
    mem[670] = 8'h00;
    mem[671] = 8'h00;
    mem[672] = 8'h00;
    mem[673] = 8'h00;
    mem[674] = 8'h00;
    mem[675] = 8'h00;
    mem[676] = 8'h00;
    mem[677] = 8'h00;
    mem[678] = 8'h00;
    mem[679] = 8'h00;
    mem[680] = 8'h00;
    mem[681] = 8'h00;
    mem[682] = 8'h00;
    mem[683] = 8'h00;
    mem[684] = 8'h00;
    mem[685] = 8'hfe;
    mem[686] = 8'hff;
    mem[687] = 8'h03;
    mem[688] = 8'hfc;
    mem[689] = 8'hff;
    mem[690] = 8'h07;
    mem[691] = 8'h00;
    mem[692] = 8'h00;
    mem[693] = 8'h00;
    mem[694] = 8'h00;
    mem[695] = 8'h00;
    mem[696] = 8'h00;
    mem[697] = 8'h00;
    mem[698] = 8'h00;
    mem[699] = 8'h00;
    mem[700] = 8'h00;
    mem[701] = 8'h00;
    mem[702] = 8'h00;
    mem[703] = 8'h00;
    mem[704] = 8'h00;
    mem[705] = 8'h00;
    mem[706] = 8'h00;
    mem[707] = 8'h00;
    mem[708] = 8'h00;
    mem[709] = 8'h00;
    mem[710] = 8'h00;
    mem[711] = 8'h00;
    mem[712] = 8'h00;
    mem[713] = 8'h00;
    mem[714] = 8'h00;
    mem[715] = 8'h00;
    mem[716] = 8'h80;
    mem[717] = 8'hff;
    mem[718] = 8'h7f;
    mem[719] = 8'h00;
    mem[720] = 8'hf0;
    mem[721] = 8'hff;
    mem[722] = 8'h1f;
    mem[723] = 8'h00;
    mem[724] = 8'h00;
    mem[725] = 8'h00;
    mem[726] = 8'h00;
    mem[727] = 8'h00;
    mem[728] = 8'h00;
    mem[729] = 8'h00;
    mem[730] = 8'h00;
    mem[731] = 8'h00;
    mem[732] = 8'h00;
    mem[733] = 8'h00;
    mem[734] = 8'h00;
    mem[735] = 8'h00;
    mem[736] = 8'h00;
    mem[737] = 8'h00;
    mem[738] = 8'h00;
    mem[739] = 8'h00;
    mem[740] = 8'h00;
    mem[741] = 8'h00;
    mem[742] = 8'h00;
    mem[743] = 8'h00;
    mem[744] = 8'h00;
    mem[745] = 8'h00;
    mem[746] = 8'h00;
    mem[747] = 8'h00;
    mem[748] = 8'h80;
    mem[749] = 8'hff;
    mem[750] = 8'h1f;
    mem[751] = 8'h00;
    mem[752] = 8'hc0;
    mem[753] = 8'hff;
    mem[754] = 8'h7f;
    mem[755] = 8'h00;
    mem[756] = 8'h00;
    mem[757] = 8'h00;
    mem[758] = 8'h00;
    mem[759] = 8'h00;
    mem[760] = 8'h00;
    mem[761] = 8'h00;
    mem[762] = 8'h00;
    mem[763] = 8'h00;
    mem[764] = 8'h00;
    mem[765] = 8'h00;
    mem[766] = 8'h00;
    mem[767] = 8'h00;
    mem[768] = 8'h00;
    mem[769] = 8'h00;
    mem[770] = 8'h00;
    mem[771] = 8'h00;
    mem[772] = 8'h00;
    mem[773] = 8'h00;
    mem[774] = 8'h00;
    mem[775] = 8'h00;
    mem[776] = 8'h00;
    mem[777] = 8'h00;
    mem[778] = 8'h00;
    mem[779] = 8'h00;
    mem[780] = 8'h80;
    mem[781] = 8'hff;
    mem[782] = 8'h07;
    mem[783] = 8'h00;
    mem[784] = 8'h00;
    mem[785] = 8'hff;
    mem[786] = 8'hff;
    mem[787] = 8'h01;
    mem[788] = 8'h00;
    mem[789] = 8'h00;
    mem[790] = 8'h00;
    mem[791] = 8'h00;
    mem[792] = 8'h00;
    mem[793] = 8'h00;
    mem[794] = 8'h00;
    mem[795] = 8'h00;
    mem[796] = 8'h00;
    mem[797] = 8'h00;
    mem[798] = 8'h00;
    mem[799] = 8'h00;
    mem[800] = 8'h00;
    mem[801] = 8'h00;
    mem[802] = 8'h00;
    mem[803] = 8'h00;
    mem[804] = 8'h00;
    mem[805] = 8'h00;
    mem[806] = 8'h00;
    mem[807] = 8'h00;
    mem[808] = 8'h00;
    mem[809] = 8'h00;
    mem[810] = 8'h00;
    mem[811] = 8'h00;
    mem[812] = 8'h00;
    mem[813] = 8'hff;
    mem[814] = 8'h01;
    mem[815] = 8'h00;
    mem[816] = 8'h00;
    mem[817] = 8'hfc;
    mem[818] = 8'hff;
    mem[819] = 8'h03;
    mem[820] = 8'h00;
    mem[821] = 8'h00;
    mem[822] = 8'h00;
    mem[823] = 8'h00;
    mem[824] = 8'h00;
    mem[825] = 8'h00;
    mem[826] = 8'h00;
    mem[827] = 8'h00;
    mem[828] = 8'h00;
    mem[829] = 8'h00;
    mem[830] = 8'h00;
    mem[831] = 8'h00;
    mem[832] = 8'h00;
    mem[833] = 8'h00;
    mem[834] = 8'h00;
    mem[835] = 8'h00;
    mem[836] = 8'h00;
    mem[837] = 8'h00;
    mem[838] = 8'h00;
    mem[839] = 8'h00;
    mem[840] = 8'h00;
    mem[841] = 8'h00;
    mem[842] = 8'h00;
    mem[843] = 8'h00;
    mem[844] = 8'h00;
    mem[845] = 8'hfe;
    mem[846] = 8'h00;
    mem[847] = 8'h00;
    mem[848] = 8'h00;
    mem[849] = 8'hf0;
    mem[850] = 8'hff;
    mem[851] = 8'h0f;
    mem[852] = 8'h00;
    mem[853] = 8'h00;
    mem[854] = 8'h00;
    mem[855] = 8'h00;
    mem[856] = 8'h00;
    mem[857] = 8'h00;
    mem[858] = 8'h00;
    mem[859] = 8'h00;
    mem[860] = 8'h00;
    mem[861] = 8'h00;
    mem[862] = 8'h00;
    mem[863] = 8'h00;
    mem[864] = 8'h00;
    mem[865] = 8'h00;
    mem[866] = 8'h00;
    mem[867] = 8'h00;
    mem[868] = 8'h00;
    mem[869] = 8'h00;
    mem[870] = 8'h00;
    mem[871] = 8'h00;
    mem[872] = 8'h00;
    mem[873] = 8'h00;
    mem[874] = 8'he0;
    mem[875] = 8'h00;
    mem[876] = 8'h00;
    mem[877] = 8'h3e;
    mem[878] = 8'h00;
    mem[879] = 8'h00;
    mem[880] = 8'h00;
    mem[881] = 8'hc0;
    mem[882] = 8'hff;
    mem[883] = 8'h3f;
    mem[884] = 8'h00;
    mem[885] = 8'h00;
    mem[886] = 8'h00;
    mem[887] = 8'h00;
    mem[888] = 8'h00;
    mem[889] = 8'h00;
    mem[890] = 8'h00;
    mem[891] = 8'h00;
    mem[892] = 8'h00;
    mem[893] = 8'h00;
    mem[894] = 8'h00;
    mem[895] = 8'h00;
    mem[896] = 8'h00;
    mem[897] = 8'h00;
    mem[898] = 8'h00;
    mem[899] = 8'h00;
    mem[900] = 8'h00;
    mem[901] = 8'h00;
    mem[902] = 8'h00;
    mem[903] = 8'h00;
    mem[904] = 8'h00;
    mem[905] = 8'h00;
    mem[906] = 8'hfc;
    mem[907] = 8'h07;
    mem[908] = 8'h00;
    mem[909] = 8'h0c;
    mem[910] = 8'h00;
    mem[911] = 8'h00;
    mem[912] = 8'h00;
    mem[913] = 8'h00;
    mem[914] = 8'hff;
    mem[915] = 8'hff;
    mem[916] = 8'h00;
    mem[917] = 8'h00;
    mem[918] = 8'h00;
    mem[919] = 8'h00;
    mem[920] = 8'h00;
    mem[921] = 8'h00;
    mem[922] = 8'h00;
    mem[923] = 8'h00;
    mem[924] = 8'h00;
    mem[925] = 8'h00;
    mem[926] = 8'h00;
    mem[927] = 8'h00;
    mem[928] = 8'h00;
    mem[929] = 8'h00;
    mem[930] = 8'h00;
    mem[931] = 8'h00;
    mem[932] = 8'h00;
    mem[933] = 8'h00;
    mem[934] = 8'h00;
    mem[935] = 8'h00;
    mem[936] = 8'h00;
    mem[937] = 8'h00;
    mem[938] = 8'hfe;
    mem[939] = 8'h0f;
    mem[940] = 8'h00;
    mem[941] = 8'h00;
    mem[942] = 8'h00;
    mem[943] = 8'h00;
    mem[944] = 8'h00;
    mem[945] = 8'h00;
    mem[946] = 8'hfc;
    mem[947] = 8'hff;
    mem[948] = 8'h03;
    mem[949] = 8'h00;
    mem[950] = 8'h00;
    mem[951] = 8'h00;
    mem[952] = 8'h00;
    mem[953] = 8'h00;
    mem[954] = 8'h00;
    mem[955] = 8'h00;
    mem[956] = 8'h00;
    mem[957] = 8'h00;
    mem[958] = 8'h00;
    mem[959] = 8'h00;
    mem[960] = 8'h00;
    mem[961] = 8'h00;
    mem[962] = 8'h00;
    mem[963] = 8'h00;
    mem[964] = 8'h00;
    mem[965] = 8'h00;
    mem[966] = 8'h00;
    mem[967] = 8'h00;
    mem[968] = 8'h00;
    mem[969] = 8'h00;
    mem[970] = 8'hff;
    mem[971] = 8'h1f;
    mem[972] = 8'h00;
    mem[973] = 8'h00;
    mem[974] = 8'h00;
    mem[975] = 8'h60;
    mem[976] = 8'h00;
    mem[977] = 8'h00;
    mem[978] = 8'hf8;
    mem[979] = 8'hff;
    mem[980] = 8'h07;
    mem[981] = 8'h00;
    mem[982] = 8'h00;
    mem[983] = 8'h00;
    mem[984] = 8'h00;
    mem[985] = 8'h00;
    mem[986] = 8'h00;
    mem[987] = 8'h00;
    mem[988] = 8'h00;
    mem[989] = 8'h00;
    mem[990] = 8'h00;
    mem[991] = 8'h00;
    mem[992] = 8'h00;
    mem[993] = 8'h00;
    mem[994] = 8'h00;
    mem[995] = 8'h00;
    mem[996] = 8'h00;
    mem[997] = 8'h00;
    mem[998] = 8'h00;
    mem[999] = 8'h00;
    mem[1000] = 8'h00;
    mem[1001] = 8'h80;
    mem[1002] = 8'hff;
    mem[1003] = 8'h3f;
    mem[1004] = 8'h00;
    mem[1005] = 8'h00;
    mem[1006] = 8'h00;
    mem[1007] = 8'hfc;
    mem[1008] = 8'h03;
    mem[1009] = 8'h00;
    mem[1010] = 8'he0;
    mem[1011] = 8'hff;
    mem[1012] = 8'h1f;
    mem[1013] = 8'h00;
    mem[1014] = 8'h00;
    mem[1015] = 8'h00;
    mem[1016] = 8'h00;
    mem[1017] = 8'h00;
    mem[1018] = 8'h00;
    mem[1019] = 8'h00;
    mem[1020] = 8'h00;
    mem[1021] = 8'h00;
    mem[1022] = 8'h00;
    mem[1023] = 8'h00;
    mem[1024] = 8'h00;
    mem[1025] = 8'h00;
    mem[1026] = 8'h00;
    mem[1027] = 8'h00;
    mem[1028] = 8'h00;
    mem[1029] = 8'h00;
    mem[1030] = 8'h00;
    mem[1031] = 8'h00;
    mem[1032] = 8'h00;
    mem[1033] = 8'hc0;
    mem[1034] = 8'h0f;
    mem[1035] = 8'h3f;
    mem[1036] = 8'h00;
    mem[1037] = 8'h00;
    mem[1038] = 8'h80;
    mem[1039] = 8'hff;
    mem[1040] = 8'h0f;
    mem[1041] = 8'h00;
    mem[1042] = 8'h80;
    mem[1043] = 8'hff;
    mem[1044] = 8'h7f;
    mem[1045] = 8'h00;
    mem[1046] = 8'h00;
    mem[1047] = 8'h00;
    mem[1048] = 8'h00;
    mem[1049] = 8'h00;
    mem[1050] = 8'h00;
    mem[1051] = 8'h00;
    mem[1052] = 8'h00;
    mem[1053] = 8'h00;
    mem[1054] = 8'h00;
    mem[1055] = 8'h00;
    mem[1056] = 8'h00;
    mem[1057] = 8'h00;
    mem[1058] = 8'h00;
    mem[1059] = 8'h00;
    mem[1060] = 8'h00;
    mem[1061] = 8'h00;
    mem[1062] = 8'h00;
    mem[1063] = 8'h00;
    mem[1064] = 8'h00;
    mem[1065] = 8'hc0;
    mem[1066] = 8'h07;
    mem[1067] = 8'h7c;
    mem[1068] = 8'h00;
    mem[1069] = 8'h00;
    mem[1070] = 8'he0;
    mem[1071] = 8'hff;
    mem[1072] = 8'h3f;
    mem[1073] = 8'h00;
    mem[1074] = 8'h00;
    mem[1075] = 8'hfe;
    mem[1076] = 8'hff;
    mem[1077] = 8'h01;
    mem[1078] = 8'h00;
    mem[1079] = 8'h00;
    mem[1080] = 8'h00;
    mem[1081] = 8'h00;
    mem[1082] = 8'h00;
    mem[1083] = 8'h00;
    mem[1084] = 8'h00;
    mem[1085] = 8'h00;
    mem[1086] = 8'h00;
    mem[1087] = 8'h00;
    mem[1088] = 8'h00;
    mem[1089] = 8'h00;
    mem[1090] = 8'h00;
    mem[1091] = 8'h00;
    mem[1092] = 8'h00;
    mem[1093] = 8'h00;
    mem[1094] = 8'h00;
    mem[1095] = 8'h00;
    mem[1096] = 8'h00;
    mem[1097] = 8'hc0;
    mem[1098] = 8'h07;
    mem[1099] = 8'h7c;
    mem[1100] = 8'h00;
    mem[1101] = 8'h00;
    mem[1102] = 8'hf8;
    mem[1103] = 8'hff;
    mem[1104] = 8'hff;
    mem[1105] = 8'h00;
    mem[1106] = 8'h00;
    mem[1107] = 8'hf8;
    mem[1108] = 8'hff;
    mem[1109] = 8'h07;
    mem[1110] = 8'h00;
    mem[1111] = 8'h00;
    mem[1112] = 8'h00;
    mem[1113] = 8'h00;
    mem[1114] = 8'h00;
    mem[1115] = 8'h00;
    mem[1116] = 8'h00;
    mem[1117] = 8'h00;
    mem[1118] = 8'h00;
    mem[1119] = 8'h00;
    mem[1120] = 8'h00;
    mem[1121] = 8'h00;
    mem[1122] = 8'h00;
    mem[1123] = 8'h00;
    mem[1124] = 8'h00;
    mem[1125] = 8'h00;
    mem[1126] = 8'h00;
    mem[1127] = 8'h00;
    mem[1128] = 8'h00;
    mem[1129] = 8'hc0;
    mem[1130] = 8'h03;
    mem[1131] = 8'h7c;
    mem[1132] = 8'h00;
    mem[1133] = 8'h00;
    mem[1134] = 8'hfe;
    mem[1135] = 8'hff;
    mem[1136] = 8'hff;
    mem[1137] = 8'h03;
    mem[1138] = 8'h00;
    mem[1139] = 8'hf0;
    mem[1140] = 8'hff;
    mem[1141] = 8'h0f;
    mem[1142] = 8'h00;
    mem[1143] = 8'h00;
    mem[1144] = 8'h00;
    mem[1145] = 8'h00;
    mem[1146] = 8'h00;
    mem[1147] = 8'h00;
    mem[1148] = 8'h00;
    mem[1149] = 8'h00;
    mem[1150] = 8'h00;
    mem[1151] = 8'h00;
    mem[1152] = 8'h00;
    mem[1153] = 8'h00;
    mem[1154] = 8'h00;
    mem[1155] = 8'h00;
    mem[1156] = 8'h00;
    mem[1157] = 8'h00;
    mem[1158] = 8'h00;
    mem[1159] = 8'h00;
    mem[1160] = 8'h00;
    mem[1161] = 8'hc0;
    mem[1162] = 8'h03;
    mem[1163] = 8'h7c;
    mem[1164] = 8'h00;
    mem[1165] = 8'h80;
    mem[1166] = 8'hff;
    mem[1167] = 8'hff;
    mem[1168] = 8'hff;
    mem[1169] = 8'h0f;
    mem[1170] = 8'h00;
    mem[1171] = 8'hc0;
    mem[1172] = 8'hff;
    mem[1173] = 8'h3f;
    mem[1174] = 8'h00;
    mem[1175] = 8'h00;
    mem[1176] = 8'h00;
    mem[1177] = 8'h00;
    mem[1178] = 8'h00;
    mem[1179] = 8'h00;
    mem[1180] = 8'h00;
    mem[1181] = 8'h00;
    mem[1182] = 8'h00;
    mem[1183] = 8'h00;
    mem[1184] = 8'h00;
    mem[1185] = 8'h00;
    mem[1186] = 8'h00;
    mem[1187] = 8'h00;
    mem[1188] = 8'h00;
    mem[1189] = 8'h00;
    mem[1190] = 8'h00;
    mem[1191] = 8'h00;
    mem[1192] = 8'h00;
    mem[1193] = 8'hf0;
    mem[1194] = 8'h07;
    mem[1195] = 8'h7c;
    mem[1196] = 8'h00;
    mem[1197] = 8'he0;
    mem[1198] = 8'hff;
    mem[1199] = 8'hff;
    mem[1200] = 8'hff;
    mem[1201] = 8'h3f;
    mem[1202] = 8'h00;
    mem[1203] = 8'h00;
    mem[1204] = 8'hff;
    mem[1205] = 8'hff;
    mem[1206] = 8'h00;
    mem[1207] = 8'h00;
    mem[1208] = 8'h00;
    mem[1209] = 8'h00;
    mem[1210] = 8'h00;
    mem[1211] = 8'h00;
    mem[1212] = 8'h00;
    mem[1213] = 8'h00;
    mem[1214] = 8'h00;
    mem[1215] = 8'h00;
    mem[1216] = 8'h00;
    mem[1217] = 8'h00;
    mem[1218] = 8'h00;
    mem[1219] = 8'h00;
    mem[1220] = 8'h00;
    mem[1221] = 8'h00;
    mem[1222] = 8'h00;
    mem[1223] = 8'h00;
    mem[1224] = 8'h00;
    mem[1225] = 8'hfc;
    mem[1226] = 8'h07;
    mem[1227] = 8'h7c;
    mem[1228] = 8'h00;
    mem[1229] = 8'hf8;
    mem[1230] = 8'hff;
    mem[1231] = 8'h8f;
    mem[1232] = 8'hff;
    mem[1233] = 8'hff;
    mem[1234] = 8'h00;
    mem[1235] = 8'h00;
    mem[1236] = 8'hfc;
    mem[1237] = 8'hff;
    mem[1238] = 8'h01;
    mem[1239] = 8'h00;
    mem[1240] = 8'h00;
    mem[1241] = 8'h00;
    mem[1242] = 8'h00;
    mem[1243] = 8'h00;
    mem[1244] = 8'h00;
    mem[1245] = 8'h00;
    mem[1246] = 8'h00;
    mem[1247] = 8'h00;
    mem[1248] = 8'h00;
    mem[1249] = 8'h00;
    mem[1250] = 8'h00;
    mem[1251] = 8'h00;
    mem[1252] = 8'h00;
    mem[1253] = 8'h00;
    mem[1254] = 8'h00;
    mem[1255] = 8'h00;
    mem[1256] = 8'h00;
    mem[1257] = 8'hfe;
    mem[1258] = 8'h0f;
    mem[1259] = 8'h3e;
    mem[1260] = 8'h00;
    mem[1261] = 8'hfe;
    mem[1262] = 8'hff;
    mem[1263] = 8'h03;
    mem[1264] = 8'hfe;
    mem[1265] = 8'hff;
    mem[1266] = 8'h03;
    mem[1267] = 8'h00;
    mem[1268] = 8'hf8;
    mem[1269] = 8'hff;
    mem[1270] = 8'h07;
    mem[1271] = 8'h00;
    mem[1272] = 8'h00;
    mem[1273] = 8'h00;
    mem[1274] = 8'h00;
    mem[1275] = 8'h00;
    mem[1276] = 8'h00;
    mem[1277] = 8'h00;
    mem[1278] = 8'h00;
    mem[1279] = 8'h00;
    mem[1280] = 8'h00;
    mem[1281] = 8'h00;
    mem[1282] = 8'h00;
    mem[1283] = 8'h00;
    mem[1284] = 8'h00;
    mem[1285] = 8'h00;
    mem[1286] = 8'h00;
    mem[1287] = 8'h00;
    mem[1288] = 8'h80;
    mem[1289] = 8'hff;
    mem[1290] = 8'hff;
    mem[1291] = 8'h3f;
    mem[1292] = 8'h80;
    mem[1293] = 8'hff;
    mem[1294] = 8'hff;
    mem[1295] = 8'h00;
    mem[1296] = 8'hf0;
    mem[1297] = 8'hff;
    mem[1298] = 8'h0f;
    mem[1299] = 8'h00;
    mem[1300] = 8'he0;
    mem[1301] = 8'hff;
    mem[1302] = 8'h1f;
    mem[1303] = 8'h00;
    mem[1304] = 8'h00;
    mem[1305] = 8'h00;
    mem[1306] = 8'h00;
    mem[1307] = 8'h00;
    mem[1308] = 8'h00;
    mem[1309] = 8'h00;
    mem[1310] = 8'h00;
    mem[1311] = 8'h00;
    mem[1312] = 8'h00;
    mem[1313] = 8'h00;
    mem[1314] = 8'h00;
    mem[1315] = 8'h00;
    mem[1316] = 8'h00;
    mem[1317] = 8'h00;
    mem[1318] = 8'h00;
    mem[1319] = 8'h00;
    mem[1320] = 8'he0;
    mem[1321] = 8'hff;
    mem[1322] = 8'hff;
    mem[1323] = 8'h1f;
    mem[1324] = 8'hc0;
    mem[1325] = 8'hff;
    mem[1326] = 8'h3f;
    mem[1327] = 8'h00;
    mem[1328] = 8'he0;
    mem[1329] = 8'hff;
    mem[1330] = 8'h3f;
    mem[1331] = 8'h00;
    mem[1332] = 8'h80;
    mem[1333] = 8'hff;
    mem[1334] = 8'h7f;
    mem[1335] = 8'h00;
    mem[1336] = 8'h00;
    mem[1337] = 8'h00;
    mem[1338] = 8'h00;
    mem[1339] = 8'h00;
    mem[1340] = 8'h00;
    mem[1341] = 8'h00;
    mem[1342] = 8'h00;
    mem[1343] = 8'h00;
    mem[1344] = 8'h00;
    mem[1345] = 8'h00;
    mem[1346] = 8'h00;
    mem[1347] = 8'h00;
    mem[1348] = 8'h00;
    mem[1349] = 8'h00;
    mem[1350] = 8'h00;
    mem[1351] = 8'h00;
    mem[1352] = 8'hf8;
    mem[1353] = 8'hff;
    mem[1354] = 8'hff;
    mem[1355] = 8'h0f;
    mem[1356] = 8'hf0;
    mem[1357] = 8'hff;
    mem[1358] = 8'h0f;
    mem[1359] = 8'h00;
    mem[1360] = 8'h80;
    mem[1361] = 8'hff;
    mem[1362] = 8'hff;
    mem[1363] = 8'h00;
    mem[1364] = 8'h00;
    mem[1365] = 8'hfe;
    mem[1366] = 8'hff;
    mem[1367] = 8'h00;
    mem[1368] = 8'h00;
    mem[1369] = 8'h00;
    mem[1370] = 8'h00;
    mem[1371] = 8'h00;
    mem[1372] = 8'h00;
    mem[1373] = 8'h00;
    mem[1374] = 8'h00;
    mem[1375] = 8'h00;
    mem[1376] = 8'h00;
    mem[1377] = 8'h00;
    mem[1378] = 8'h00;
    mem[1379] = 8'h00;
    mem[1380] = 8'h00;
    mem[1381] = 8'h00;
    mem[1382] = 8'h00;
    mem[1383] = 8'h00;
    mem[1384] = 8'hfc;
    mem[1385] = 8'hff;
    mem[1386] = 8'hfc;
    mem[1387] = 8'h07;
    mem[1388] = 8'hfc;
    mem[1389] = 8'hff;
    mem[1390] = 8'h03;
    mem[1391] = 8'h00;
    mem[1392] = 8'h00;
    mem[1393] = 8'hfe;
    mem[1394] = 8'hff;
    mem[1395] = 8'h01;
    mem[1396] = 8'h00;
    mem[1397] = 8'hf8;
    mem[1398] = 8'hff;
    mem[1399] = 8'h03;
    mem[1400] = 8'h00;
    mem[1401] = 8'h00;
    mem[1402] = 8'h00;
    mem[1403] = 8'h00;
    mem[1404] = 8'h00;
    mem[1405] = 8'h00;
    mem[1406] = 8'h00;
    mem[1407] = 8'h00;
    mem[1408] = 8'h00;
    mem[1409] = 8'h00;
    mem[1410] = 8'h00;
    mem[1411] = 8'h00;
    mem[1412] = 8'h00;
    mem[1413] = 8'h00;
    mem[1414] = 8'h00;
    mem[1415] = 8'h00;
    mem[1416] = 8'hff;
    mem[1417] = 8'h7f;
    mem[1418] = 8'he0;
    mem[1419] = 8'h00;
    mem[1420] = 8'hff;
    mem[1421] = 8'hff;
    mem[1422] = 8'h00;
    mem[1423] = 8'h00;
    mem[1424] = 8'h00;
    mem[1425] = 8'hf8;
    mem[1426] = 8'hff;
    mem[1427] = 8'h07;
    mem[1428] = 8'h00;
    mem[1429] = 8'hf0;
    mem[1430] = 8'hff;
    mem[1431] = 8'h0f;
    mem[1432] = 8'h00;
    mem[1433] = 8'h00;
    mem[1434] = 8'h00;
    mem[1435] = 8'h00;
    mem[1436] = 8'h00;
    mem[1437] = 8'h00;
    mem[1438] = 8'h00;
    mem[1439] = 8'h00;
    mem[1440] = 8'h00;
    mem[1441] = 8'h00;
    mem[1442] = 8'h00;
    mem[1443] = 8'h00;
    mem[1444] = 8'h00;
    mem[1445] = 8'h00;
    mem[1446] = 8'h00;
    mem[1447] = 8'hc0;
    mem[1448] = 8'hff;
    mem[1449] = 8'h1f;
    mem[1450] = 8'h00;
    mem[1451] = 8'hc0;
    mem[1452] = 8'hff;
    mem[1453] = 8'h3f;
    mem[1454] = 8'h00;
    mem[1455] = 8'h20;
    mem[1456] = 8'h00;
    mem[1457] = 8'he0;
    mem[1458] = 8'hff;
    mem[1459] = 8'h1f;
    mem[1460] = 8'h00;
    mem[1461] = 8'hc0;
    mem[1462] = 8'hff;
    mem[1463] = 8'h1f;
    mem[1464] = 8'h00;
    mem[1465] = 8'h00;
    mem[1466] = 8'h00;
    mem[1467] = 8'h00;
    mem[1468] = 8'h00;
    mem[1469] = 8'h00;
    mem[1470] = 8'h00;
    mem[1471] = 8'h00;
    mem[1472] = 8'h00;
    mem[1473] = 8'h00;
    mem[1474] = 8'h00;
    mem[1475] = 8'h00;
    mem[1476] = 8'h00;
    mem[1477] = 8'h00;
    mem[1478] = 8'h00;
    mem[1479] = 8'he0;
    mem[1480] = 8'hff;
    mem[1481] = 8'h0f;
    mem[1482] = 8'h00;
    mem[1483] = 8'he0;
    mem[1484] = 8'hff;
    mem[1485] = 8'h0f;
    mem[1486] = 8'h00;
    mem[1487] = 8'hfc;
    mem[1488] = 8'h03;
    mem[1489] = 8'h80;
    mem[1490] = 8'hff;
    mem[1491] = 8'h7f;
    mem[1492] = 8'h00;
    mem[1493] = 8'h00;
    mem[1494] = 8'hff;
    mem[1495] = 8'h7f;
    mem[1496] = 8'h00;
    mem[1497] = 8'h00;
    mem[1498] = 8'h00;
    mem[1499] = 8'h00;
    mem[1500] = 8'h00;
    mem[1501] = 8'h00;
    mem[1502] = 8'h00;
    mem[1503] = 8'h00;
    mem[1504] = 8'h00;
    mem[1505] = 8'h00;
    mem[1506] = 8'h00;
    mem[1507] = 8'h00;
    mem[1508] = 8'h00;
    mem[1509] = 8'h00;
    mem[1510] = 8'h00;
    mem[1511] = 8'hf8;
    mem[1512] = 8'hff;
    mem[1513] = 8'h03;
    mem[1514] = 8'h00;
    mem[1515] = 8'hf8;
    mem[1516] = 8'hff;
    mem[1517] = 8'h07;
    mem[1518] = 8'h00;
    mem[1519] = 8'hff;
    mem[1520] = 8'h07;
    mem[1521] = 8'h00;
    mem[1522] = 8'hfe;
    mem[1523] = 8'hff;
    mem[1524] = 8'h01;
    mem[1525] = 8'h00;
    mem[1526] = 8'hfe;
    mem[1527] = 8'hff;
    mem[1528] = 8'h00;
    mem[1529] = 8'h00;
    mem[1530] = 8'h00;
    mem[1531] = 8'h00;
    mem[1532] = 8'h00;
    mem[1533] = 8'h00;
    mem[1534] = 8'h00;
    mem[1535] = 8'h00;
    mem[1536] = 8'h00;
    mem[1537] = 8'h00;
    mem[1538] = 8'h00;
    mem[1539] = 8'h00;
    mem[1540] = 8'h00;
    mem[1541] = 8'h00;
    mem[1542] = 8'h00;
    mem[1543] = 8'hfc;
    mem[1544] = 8'hff;
    mem[1545] = 8'h00;
    mem[1546] = 8'h00;
    mem[1547] = 8'hfe;
    mem[1548] = 8'hff;
    mem[1549] = 8'h01;
    mem[1550] = 8'h80;
    mem[1551] = 8'hff;
    mem[1552] = 8'h0f;
    mem[1553] = 8'h00;
    mem[1554] = 8'hf8;
    mem[1555] = 8'hff;
    mem[1556] = 8'h03;
    mem[1557] = 8'h00;
    mem[1558] = 8'hf8;
    mem[1559] = 8'hff;
    mem[1560] = 8'h03;
    mem[1561] = 8'h00;
    mem[1562] = 8'h00;
    mem[1563] = 8'h00;
    mem[1564] = 8'h00;
    mem[1565] = 8'h00;
    mem[1566] = 8'h00;
    mem[1567] = 8'h00;
    mem[1568] = 8'h00;
    mem[1569] = 8'h00;
    mem[1570] = 8'h00;
    mem[1571] = 8'h00;
    mem[1572] = 8'h00;
    mem[1573] = 8'h00;
    mem[1574] = 8'h00;
    mem[1575] = 8'hff;
    mem[1576] = 8'h7f;
    mem[1577] = 8'h00;
    mem[1578] = 8'h80;
    mem[1579] = 8'hff;
    mem[1580] = 8'h7f;
    mem[1581] = 8'h00;
    mem[1582] = 8'hc0;
    mem[1583] = 8'h07;
    mem[1584] = 8'h1e;
    mem[1585] = 8'h00;
    mem[1586] = 8'hf0;
    mem[1587] = 8'hff;
    mem[1588] = 8'h0f;
    mem[1589] = 8'h00;
    mem[1590] = 8'he0;
    mem[1591] = 8'hff;
    mem[1592] = 8'h0f;
    mem[1593] = 8'h00;
    mem[1594] = 8'h00;
    mem[1595] = 8'h00;
    mem[1596] = 8'h00;
    mem[1597] = 8'h00;
    mem[1598] = 8'h00;
    mem[1599] = 8'h00;
    mem[1600] = 8'h00;
    mem[1601] = 8'h00;
    mem[1602] = 8'h00;
    mem[1603] = 8'h00;
    mem[1604] = 8'h00;
    mem[1605] = 8'h00;
    mem[1606] = 8'hc0;
    mem[1607] = 8'hff;
    mem[1608] = 8'h1f;
    mem[1609] = 8'h00;
    mem[1610] = 8'hc0;
    mem[1611] = 8'hff;
    mem[1612] = 8'h1f;
    mem[1613] = 8'h00;
    mem[1614] = 8'he0;
    mem[1615] = 8'hf9;
    mem[1616] = 8'h1c;
    mem[1617] = 8'h00;
    mem[1618] = 8'hc0;
    mem[1619] = 8'hff;
    mem[1620] = 8'h3f;
    mem[1621] = 8'h00;
    mem[1622] = 8'hc0;
    mem[1623] = 8'hff;
    mem[1624] = 8'h1f;
    mem[1625] = 8'h00;
    mem[1626] = 8'h00;
    mem[1627] = 8'h00;
    mem[1628] = 8'h00;
    mem[1629] = 8'h00;
    mem[1630] = 8'h00;
    mem[1631] = 8'h00;
    mem[1632] = 8'h00;
    mem[1633] = 8'h00;
    mem[1634] = 8'h00;
    mem[1635] = 8'h00;
    mem[1636] = 8'h00;
    mem[1637] = 8'h00;
    mem[1638] = 8'he0;
    mem[1639] = 8'hff;
    mem[1640] = 8'h07;
    mem[1641] = 8'h00;
    mem[1642] = 8'hf0;
    mem[1643] = 8'hff;
    mem[1644] = 8'h07;
    mem[1645] = 8'h00;
    mem[1646] = 8'hf8;
    mem[1647] = 8'hf9;
    mem[1648] = 8'h39;
    mem[1649] = 8'h00;
    mem[1650] = 8'h00;
    mem[1651] = 8'hff;
    mem[1652] = 8'hff;
    mem[1653] = 8'h00;
    mem[1654] = 8'h00;
    mem[1655] = 8'hff;
    mem[1656] = 8'h7f;
    mem[1657] = 8'h00;
    mem[1658] = 8'h00;
    mem[1659] = 8'h00;
    mem[1660] = 8'h00;
    mem[1661] = 8'h00;
    mem[1662] = 8'h00;
    mem[1663] = 8'h00;
    mem[1664] = 8'h00;
    mem[1665] = 8'h00;
    mem[1666] = 8'h00;
    mem[1667] = 8'h00;
    mem[1668] = 8'h00;
    mem[1669] = 8'h00;
    mem[1670] = 8'hf8;
    mem[1671] = 8'hff;
    mem[1672] = 8'h01;
    mem[1673] = 8'h00;
    mem[1674] = 8'hfc;
    mem[1675] = 8'hff;
    mem[1676] = 8'h03;
    mem[1677] = 8'h00;
    mem[1678] = 8'hfc;
    mem[1679] = 8'hfc;
    mem[1680] = 8'h39;
    mem[1681] = 8'h00;
    mem[1682] = 8'h00;
    mem[1683] = 8'hfc;
    mem[1684] = 8'hff;
    mem[1685] = 8'h01;
    mem[1686] = 8'h00;
    mem[1687] = 8'hfc;
    mem[1688] = 8'hff;
    mem[1689] = 8'h00;
    mem[1690] = 8'h00;
    mem[1691] = 8'h00;
    mem[1692] = 8'h00;
    mem[1693] = 8'h00;
    mem[1694] = 8'h00;
    mem[1695] = 8'h00;
    mem[1696] = 8'h00;
    mem[1697] = 8'h00;
    mem[1698] = 8'h00;
    mem[1699] = 8'h00;
    mem[1700] = 8'h00;
    mem[1701] = 8'h00;
    mem[1702] = 8'hfc;
    mem[1703] = 8'hff;
    mem[1704] = 8'h00;
    mem[1705] = 8'h00;
    mem[1706] = 8'hfe;
    mem[1707] = 8'hff;
    mem[1708] = 8'h00;
    mem[1709] = 8'h00;
    mem[1710] = 8'hff;
    mem[1711] = 8'h9c;
    mem[1712] = 8'h3b;
    mem[1713] = 8'h00;
    mem[1714] = 8'h00;
    mem[1715] = 8'hf8;
    mem[1716] = 8'hff;
    mem[1717] = 8'h07;
    mem[1718] = 8'h00;
    mem[1719] = 8'hf8;
    mem[1720] = 8'hff;
    mem[1721] = 8'h03;
    mem[1722] = 8'h00;
    mem[1723] = 8'h00;
    mem[1724] = 8'h00;
    mem[1725] = 8'h00;
    mem[1726] = 8'h00;
    mem[1727] = 8'h00;
    mem[1728] = 8'h00;
    mem[1729] = 8'h00;
    mem[1730] = 8'h00;
    mem[1731] = 8'h00;
    mem[1732] = 8'h00;
    mem[1733] = 8'h00;
    mem[1734] = 8'hff;
    mem[1735] = 8'h3f;
    mem[1736] = 8'h00;
    mem[1737] = 8'h80;
    mem[1738] = 8'hff;
    mem[1739] = 8'h3f;
    mem[1740] = 8'h00;
    mem[1741] = 8'hc0;
    mem[1742] = 8'hef;
    mem[1743] = 8'hdc;
    mem[1744] = 8'h3b;
    mem[1745] = 8'h00;
    mem[1746] = 8'h00;
    mem[1747] = 8'he0;
    mem[1748] = 8'hff;
    mem[1749] = 8'h1f;
    mem[1750] = 8'h00;
    mem[1751] = 8'he0;
    mem[1752] = 8'hff;
    mem[1753] = 8'h07;
    mem[1754] = 8'h00;
    mem[1755] = 8'h00;
    mem[1756] = 8'h00;
    mem[1757] = 8'h00;
    mem[1758] = 8'h00;
    mem[1759] = 8'h00;
    mem[1760] = 8'h00;
    mem[1761] = 8'h00;
    mem[1762] = 8'h00;
    mem[1763] = 8'h00;
    mem[1764] = 8'h00;
    mem[1765] = 8'h80;
    mem[1766] = 8'hff;
    mem[1767] = 8'h1f;
    mem[1768] = 8'h00;
    mem[1769] = 8'he0;
    mem[1770] = 8'hff;
    mem[1771] = 8'h1f;
    mem[1772] = 8'h00;
    mem[1773] = 8'hf0;
    mem[1774] = 8'he7;
    mem[1775] = 8'hfc;
    mem[1776] = 8'h39;
    mem[1777] = 8'h00;
    mem[1778] = 8'h00;
    mem[1779] = 8'h80;
    mem[1780] = 8'hff;
    mem[1781] = 8'h3f;
    mem[1782] = 8'h00;
    mem[1783] = 8'h80;
    mem[1784] = 8'hff;
    mem[1785] = 8'h1f;
    mem[1786] = 8'h00;
    mem[1787] = 8'h00;
    mem[1788] = 8'h00;
    mem[1789] = 8'h00;
    mem[1790] = 8'h00;
    mem[1791] = 8'h00;
    mem[1792] = 8'h00;
    mem[1793] = 8'h00;
    mem[1794] = 8'h00;
    mem[1795] = 8'h00;
    mem[1796] = 8'h00;
    mem[1797] = 8'he0;
    mem[1798] = 8'hff;
    mem[1799] = 8'h07;
    mem[1800] = 8'h00;
    mem[1801] = 8'hf0;
    mem[1802] = 8'hff;
    mem[1803] = 8'h07;
    mem[1804] = 8'h00;
    mem[1805] = 8'hf8;
    mem[1806] = 8'hc1;
    mem[1807] = 8'hf9;
    mem[1808] = 8'h3d;
    mem[1809] = 8'h00;
    mem[1810] = 8'h00;
    mem[1811] = 8'h00;
    mem[1812] = 8'hff;
    mem[1813] = 8'hff;
    mem[1814] = 8'h00;
    mem[1815] = 8'h00;
    mem[1816] = 8'hff;
    mem[1817] = 8'h3f;
    mem[1818] = 8'h00;
    mem[1819] = 8'h00;
    mem[1820] = 8'h00;
    mem[1821] = 8'h00;
    mem[1822] = 8'h00;
    mem[1823] = 8'h00;
    mem[1824] = 8'h00;
    mem[1825] = 8'h00;
    mem[1826] = 8'h00;
    mem[1827] = 8'h00;
    mem[1828] = 8'h00;
    mem[1829] = 8'hf0;
    mem[1830] = 8'hff;
    mem[1831] = 8'h01;
    mem[1832] = 8'h00;
    mem[1833] = 8'hfc;
    mem[1834] = 8'hff;
    mem[1835] = 8'h01;
    mem[1836] = 8'h00;
    mem[1837] = 8'h7e;
    mem[1838] = 8'hc0;
    mem[1839] = 8'hf3;
    mem[1840] = 8'h1c;
    mem[1841] = 8'h00;
    mem[1842] = 8'h00;
    mem[1843] = 8'h00;
    mem[1844] = 8'hfc;
    mem[1845] = 8'hff;
    mem[1846] = 8'h03;
    mem[1847] = 8'h00;
    mem[1848] = 8'hfc;
    mem[1849] = 8'hff;
    mem[1850] = 8'h00;
    mem[1851] = 8'h00;
    mem[1852] = 8'h00;
    mem[1853] = 8'h00;
    mem[1854] = 8'h00;
    mem[1855] = 8'h00;
    mem[1856] = 8'h00;
    mem[1857] = 8'h00;
    mem[1858] = 8'h00;
    mem[1859] = 8'h00;
    mem[1860] = 8'h00;
    mem[1861] = 8'hfc;
    mem[1862] = 8'hff;
    mem[1863] = 8'h00;
    mem[1864] = 8'h00;
    mem[1865] = 8'hff;
    mem[1866] = 8'h7f;
    mem[1867] = 8'h00;
    mem[1868] = 8'h80;
    mem[1869] = 8'h1f;
    mem[1870] = 8'h80;
    mem[1871] = 8'h07;
    mem[1872] = 8'h1e;
    mem[1873] = 8'h00;
    mem[1874] = 8'hc0;
    mem[1875] = 8'h1f;
    mem[1876] = 8'hf0;
    mem[1877] = 8'hff;
    mem[1878] = 8'h07;
    mem[1879] = 8'h00;
    mem[1880] = 8'hf8;
    mem[1881] = 8'hff;
    mem[1882] = 8'h01;
    mem[1883] = 8'h00;
    mem[1884] = 8'h00;
    mem[1885] = 8'h00;
    mem[1886] = 8'h00;
    mem[1887] = 8'h00;
    mem[1888] = 8'h00;
    mem[1889] = 8'h00;
    mem[1890] = 8'h00;
    mem[1891] = 8'h00;
    mem[1892] = 8'h00;
    mem[1893] = 8'hfe;
    mem[1894] = 8'h3f;
    mem[1895] = 8'h00;
    mem[1896] = 8'h80;
    mem[1897] = 8'hff;
    mem[1898] = 8'h3f;
    mem[1899] = 8'h00;
    mem[1900] = 8'he0;
    mem[1901] = 8'h07;
    mem[1902] = 8'h80;
    mem[1903] = 8'hff;
    mem[1904] = 8'h0f;
    mem[1905] = 8'h00;
    mem[1906] = 8'he0;
    mem[1907] = 8'h7f;
    mem[1908] = 8'hc0;
    mem[1909] = 8'hff;
    mem[1910] = 8'h1f;
    mem[1911] = 8'h00;
    mem[1912] = 8'he0;
    mem[1913] = 8'hff;
    mem[1914] = 8'h07;
    mem[1915] = 8'h00;
    mem[1916] = 8'h00;
    mem[1917] = 8'h00;
    mem[1918] = 8'h00;
    mem[1919] = 8'h00;
    mem[1920] = 8'h00;
    mem[1921] = 8'h00;
    mem[1922] = 8'h00;
    mem[1923] = 8'h00;
    mem[1924] = 8'h00;
    mem[1925] = 8'hff;
    mem[1926] = 8'h1f;
    mem[1927] = 8'h00;
    mem[1928] = 8'he0;
    mem[1929] = 8'hff;
    mem[1930] = 8'h0f;
    mem[1931] = 8'h00;
    mem[1932] = 8'hf3;
    mem[1933] = 8'h03;
    mem[1934] = 8'h80;
    mem[1935] = 8'hff;
    mem[1936] = 8'h0f;
    mem[1937] = 8'h00;
    mem[1938] = 8'hf8;
    mem[1939] = 8'hff;
    mem[1940] = 8'h80;
    mem[1941] = 8'hff;
    mem[1942] = 8'h3f;
    mem[1943] = 8'h00;
    mem[1944] = 8'h80;
    mem[1945] = 8'hff;
    mem[1946] = 8'h0f;
    mem[1947] = 8'h00;
    mem[1948] = 8'h00;
    mem[1949] = 8'h00;
    mem[1950] = 8'h00;
    mem[1951] = 8'h00;
    mem[1952] = 8'h00;
    mem[1953] = 8'h00;
    mem[1954] = 8'h00;
    mem[1955] = 8'h00;
    mem[1956] = 8'hc0;
    mem[1957] = 8'hff;
    mem[1958] = 8'h07;
    mem[1959] = 8'h00;
    mem[1960] = 8'hf8;
    mem[1961] = 8'hff;
    mem[1962] = 8'h03;
    mem[1963] = 8'he0;
    mem[1964] = 8'hff;
    mem[1965] = 8'h00;
    mem[1966] = 8'hc0;
    mem[1967] = 8'hff;
    mem[1968] = 8'h0f;
    mem[1969] = 8'h00;
    mem[1970] = 8'hf8;
    mem[1971] = 8'hff;
    mem[1972] = 8'h01;
    mem[1973] = 8'hfe;
    mem[1974] = 8'hff;
    mem[1975] = 8'h00;
    mem[1976] = 8'h00;
    mem[1977] = 8'hff;
    mem[1978] = 8'h1f;
    mem[1979] = 8'h00;
    mem[1980] = 8'h00;
    mem[1981] = 8'h00;
    mem[1982] = 8'h00;
    mem[1983] = 8'h00;
    mem[1984] = 8'h00;
    mem[1985] = 8'h00;
    mem[1986] = 8'h00;
    mem[1987] = 8'h00;
    mem[1988] = 8'he0;
    mem[1989] = 8'hff;
    mem[1990] = 8'h03;
    mem[1991] = 8'h00;
    mem[1992] = 8'hfc;
    mem[1993] = 8'hff;
    mem[1994] = 8'h00;
    mem[1995] = 8'hf8;
    mem[1996] = 8'h7f;
    mem[1997] = 8'h00;
    mem[1998] = 8'hf0;
    mem[1999] = 8'h73;
    mem[2000] = 8'h0e;
    mem[2001] = 8'h00;
    mem[2002] = 8'hfc;
    mem[2003] = 8'hfd;
    mem[2004] = 8'h01;
    mem[2005] = 8'hf8;
    mem[2006] = 8'hff;
    mem[2007] = 8'h03;
    mem[2008] = 8'h00;
    mem[2009] = 8'hfc;
    mem[2010] = 8'h3f;
    mem[2011] = 8'h00;
    mem[2012] = 8'h00;
    mem[2013] = 8'h00;
    mem[2014] = 8'h00;
    mem[2015] = 8'h00;
    mem[2016] = 8'h00;
    mem[2017] = 8'h00;
    mem[2018] = 8'h00;
    mem[2019] = 8'h00;
    mem[2020] = 8'hf0;
    mem[2021] = 8'hff;
    mem[2022] = 8'h00;
    mem[2023] = 8'h00;
    mem[2024] = 8'hff;
    mem[2025] = 8'h7f;
    mem[2026] = 8'h00;
    mem[2027] = 8'hfc;
    mem[2028] = 8'hfc;
    mem[2029] = 8'h00;
    mem[2030] = 8'hfc;
    mem[2031] = 8'h73;
    mem[2032] = 8'h0e;
    mem[2033] = 8'h00;
    mem[2034] = 8'h7c;
    mem[2035] = 8'hf0;
    mem[2036] = 8'h03;
    mem[2037] = 8'he0;
    mem[2038] = 8'hff;
    mem[2039] = 8'h07;
    mem[2040] = 8'h00;
    mem[2041] = 8'hf8;
    mem[2042] = 8'h7f;
    mem[2043] = 8'h00;
    mem[2044] = 8'h00;
    mem[2045] = 8'h00;
    mem[2046] = 8'h00;
    mem[2047] = 8'h00;
    mem[2048] = 8'h00;
    mem[2049] = 8'h00;
    mem[2050] = 8'h00;
    mem[2051] = 8'h00;
    mem[2052] = 8'hf8;
    mem[2053] = 8'h7f;
    mem[2054] = 8'h00;
    mem[2055] = 8'h80;
    mem[2056] = 8'hff;
    mem[2057] = 8'h1f;
    mem[2058] = 8'h00;
    mem[2059] = 8'h3c;
    mem[2060] = 8'hf0;
    mem[2061] = 8'h00;
    mem[2062] = 8'hff;
    mem[2063] = 8'h73;
    mem[2064] = 8'h0e;
    mem[2065] = 8'h00;
    mem[2066] = 8'h3e;
    mem[2067] = 8'he0;
    mem[2068] = 8'h03;
    mem[2069] = 8'hc0;
    mem[2070] = 8'hff;
    mem[2071] = 8'h1f;
    mem[2072] = 8'h00;
    mem[2073] = 8'he0;
    mem[2074] = 8'hff;
    mem[2075] = 8'h00;
    mem[2076] = 8'h00;
    mem[2077] = 8'h00;
    mem[2078] = 8'h00;
    mem[2079] = 8'h00;
    mem[2080] = 8'h00;
    mem[2081] = 8'h00;
    mem[2082] = 8'h00;
    mem[2083] = 8'h00;
    mem[2084] = 8'hf8;
    mem[2085] = 8'h1f;
    mem[2086] = 8'h00;
    mem[2087] = 8'he0;
    mem[2088] = 8'hff;
    mem[2089] = 8'h07;
    mem[2090] = 8'h00;
    mem[2091] = 8'h9e;
    mem[2092] = 8'he7;
    mem[2093] = 8'h81;
    mem[2094] = 8'h9f;
    mem[2095] = 8'h73;
    mem[2096] = 8'h0e;
    mem[2097] = 8'h00;
    mem[2098] = 8'h3e;
    mem[2099] = 8'hc0;
    mem[2100] = 8'h03;
    mem[2101] = 8'h00;
    mem[2102] = 8'hff;
    mem[2103] = 8'h3f;
    mem[2104] = 8'h00;
    mem[2105] = 8'hc0;
    mem[2106] = 8'hff;
    mem[2107] = 8'h01;
    mem[2108] = 8'h00;
    mem[2109] = 8'h00;
    mem[2110] = 8'h00;
    mem[2111] = 8'h00;
    mem[2112] = 8'h00;
    mem[2113] = 8'h00;
    mem[2114] = 8'h00;
    mem[2115] = 8'h00;
    mem[2116] = 8'hf8;
    mem[2117] = 8'h0f;
    mem[2118] = 8'h00;
    mem[2119] = 8'hf0;
    mem[2120] = 8'hff;
    mem[2121] = 8'h03;
    mem[2122] = 8'h00;
    mem[2123] = 8'hcf;
    mem[2124] = 8'hcf;
    mem[2125] = 8'he1;
    mem[2126] = 8'h87;
    mem[2127] = 8'h73;
    mem[2128] = 8'h0e;
    mem[2129] = 8'h00;
    mem[2130] = 8'h3e;
    mem[2131] = 8'hc0;
    mem[2132] = 8'h03;
    mem[2133] = 8'h00;
    mem[2134] = 8'hfc;
    mem[2135] = 8'hff;
    mem[2136] = 8'h00;
    mem[2137] = 8'h80;
    mem[2138] = 8'hff;
    mem[2139] = 8'h01;
    mem[2140] = 8'h00;
    mem[2141] = 8'h00;
    mem[2142] = 8'h00;
    mem[2143] = 8'h00;
    mem[2144] = 8'h00;
    mem[2145] = 8'h00;
    mem[2146] = 8'h00;
    mem[2147] = 8'h00;
    mem[2148] = 8'hfc;
    mem[2149] = 8'h07;
    mem[2150] = 8'h00;
    mem[2151] = 8'hfc;
    mem[2152] = 8'hff;
    mem[2153] = 8'h00;
    mem[2154] = 8'h80;
    mem[2155] = 8'hef;
    mem[2156] = 8'hdf;
    mem[2157] = 8'hf9;
    mem[2158] = 8'h81;
    mem[2159] = 8'hff;
    mem[2160] = 8'h0f;
    mem[2161] = 8'h00;
    mem[2162] = 8'h3e;
    mem[2163] = 8'hc0;
    mem[2164] = 8'h07;
    mem[2165] = 8'h00;
    mem[2166] = 8'hf8;
    mem[2167] = 8'hff;
    mem[2168] = 8'h01;
    mem[2169] = 8'h00;
    mem[2170] = 8'hfe;
    mem[2171] = 8'h01;
    mem[2172] = 8'h00;
    mem[2173] = 8'h00;
    mem[2174] = 8'h00;
    mem[2175] = 8'h00;
    mem[2176] = 8'h00;
    mem[2177] = 8'h00;
    mem[2178] = 8'h00;
    mem[2179] = 8'h00;
    mem[2180] = 8'hfc;
    mem[2181] = 8'h03;
    mem[2182] = 8'h00;
    mem[2183] = 8'hfe;
    mem[2184] = 8'h7f;
    mem[2185] = 8'h00;
    mem[2186] = 8'he0;
    mem[2187] = 8'hef;
    mem[2188] = 8'hdc;
    mem[2189] = 8'h7f;
    mem[2190] = 8'h80;
    mem[2191] = 8'hff;
    mem[2192] = 8'h0f;
    mem[2193] = 8'h00;
    mem[2194] = 8'h3e;
    mem[2195] = 8'he0;
    mem[2196] = 8'h0f;
    mem[2197] = 8'h00;
    mem[2198] = 8'he0;
    mem[2199] = 8'hff;
    mem[2200] = 8'h07;
    mem[2201] = 8'h00;
    mem[2202] = 8'hfe;
    mem[2203] = 8'h01;
    mem[2204] = 8'h00;
    mem[2205] = 8'h00;
    mem[2206] = 8'h00;
    mem[2207] = 8'h00;
    mem[2208] = 8'h00;
    mem[2209] = 8'h00;
    mem[2210] = 8'h00;
    mem[2211] = 8'h00;
    mem[2212] = 8'hfc;
    mem[2213] = 8'h03;
    mem[2214] = 8'h80;
    mem[2215] = 8'hff;
    mem[2216] = 8'h1f;
    mem[2217] = 8'h00;
    mem[2218] = 8'hf0;
    mem[2219] = 8'hef;
    mem[2220] = 8'hdc;
    mem[2221] = 8'h3f;
    mem[2222] = 8'h80;
    mem[2223] = 8'hff;
    mem[2224] = 8'h0f;
    mem[2225] = 8'h00;
    mem[2226] = 8'h7c;
    mem[2227] = 8'hf0;
    mem[2228] = 8'h3f;
    mem[2229] = 8'h00;
    mem[2230] = 8'h80;
    mem[2231] = 8'hff;
    mem[2232] = 8'h0f;
    mem[2233] = 8'h00;
    mem[2234] = 8'hfc;
    mem[2235] = 8'h01;
    mem[2236] = 8'h00;
    mem[2237] = 8'h00;
    mem[2238] = 8'h00;
    mem[2239] = 8'h00;
    mem[2240] = 8'h00;
    mem[2241] = 8'h00;
    mem[2242] = 8'h00;
    mem[2243] = 8'h00;
    mem[2244] = 8'hfc;
    mem[2245] = 8'h03;
    mem[2246] = 8'hc0;
    mem[2247] = 8'hff;
    mem[2248] = 8'h07;
    mem[2249] = 8'h00;
    mem[2250] = 8'hfc;
    mem[2251] = 8'hee;
    mem[2252] = 8'hdf;
    mem[2253] = 8'h0f;
    mem[2254] = 8'h00;
    mem[2255] = 8'h9c;
    mem[2256] = 8'h03;
    mem[2257] = 8'h00;
    mem[2258] = 8'hfc;
    mem[2259] = 8'hfd;
    mem[2260] = 8'hff;
    mem[2261] = 8'h00;
    mem[2262] = 8'h00;
    mem[2263] = 8'hff;
    mem[2264] = 8'h1f;
    mem[2265] = 8'h00;
    mem[2266] = 8'hfc;
    mem[2267] = 8'h01;
    mem[2268] = 8'h00;
    mem[2269] = 8'h00;
    mem[2270] = 8'h00;
    mem[2271] = 8'h00;
    mem[2272] = 8'h00;
    mem[2273] = 8'h00;
    mem[2274] = 8'h00;
    mem[2275] = 8'h00;
    mem[2276] = 8'hfc;
    mem[2277] = 8'h01;
    mem[2278] = 8'he0;
    mem[2279] = 8'hff;
    mem[2280] = 8'h03;
    mem[2281] = 8'h00;
    mem[2282] = 8'h3e;
    mem[2283] = 8'hce;
    mem[2284] = 8'hcf;
    mem[2285] = 8'h03;
    mem[2286] = 8'h00;
    mem[2287] = 8'hfc;
    mem[2288] = 8'h03;
    mem[2289] = 8'h00;
    mem[2290] = 8'hf8;
    mem[2291] = 8'hff;
    mem[2292] = 8'hff;
    mem[2293] = 8'h01;
    mem[2294] = 8'h00;
    mem[2295] = 8'hfc;
    mem[2296] = 8'h3f;
    mem[2297] = 8'h00;
    mem[2298] = 8'hfc;
    mem[2299] = 8'h03;
    mem[2300] = 8'h00;
    mem[2301] = 8'h00;
    mem[2302] = 8'h00;
    mem[2303] = 8'h00;
    mem[2304] = 8'h00;
    mem[2305] = 8'h00;
    mem[2306] = 8'h00;
    mem[2307] = 8'h00;
    mem[2308] = 8'hfc;
    mem[2309] = 8'h01;
    mem[2310] = 8'hf0;
    mem[2311] = 8'hff;
    mem[2312] = 8'h00;
    mem[2313] = 8'h80;
    mem[2314] = 8'h1f;
    mem[2315] = 8'h9e;
    mem[2316] = 8'he7;
    mem[2317] = 8'h01;
    mem[2318] = 8'h00;
    mem[2319] = 8'hfc;
    mem[2320] = 8'h03;
    mem[2321] = 8'h00;
    mem[2322] = 8'hf8;
    mem[2323] = 8'hff;
    mem[2324] = 8'hff;
    mem[2325] = 8'h07;
    mem[2326] = 8'h00;
    mem[2327] = 8'hf8;
    mem[2328] = 8'hff;
    mem[2329] = 8'h00;
    mem[2330] = 8'hfc;
    mem[2331] = 8'h03;
    mem[2332] = 8'h00;
    mem[2333] = 8'h00;
    mem[2334] = 8'h00;
    mem[2335] = 8'h00;
    mem[2336] = 8'h00;
    mem[2337] = 8'h00;
    mem[2338] = 8'h00;
    mem[2339] = 8'h00;
    mem[2340] = 8'hfc;
    mem[2341] = 8'h01;
    mem[2342] = 8'hf8;
    mem[2343] = 8'h7f;
    mem[2344] = 8'h00;
    mem[2345] = 8'hc0;
    mem[2346] = 8'h07;
    mem[2347] = 8'h3c;
    mem[2348] = 8'hf0;
    mem[2349] = 8'h00;
    mem[2350] = 8'h00;
    mem[2351] = 8'hfc;
    mem[2352] = 8'h03;
    mem[2353] = 8'h00;
    mem[2354] = 8'he0;
    mem[2355] = 8'hff;
    mem[2356] = 8'hff;
    mem[2357] = 8'h0f;
    mem[2358] = 8'h00;
    mem[2359] = 8'he0;
    mem[2360] = 8'hff;
    mem[2361] = 8'h00;
    mem[2362] = 8'hfc;
    mem[2363] = 8'h03;
    mem[2364] = 8'h00;
    mem[2365] = 8'h00;
    mem[2366] = 8'h00;
    mem[2367] = 8'h00;
    mem[2368] = 8'h00;
    mem[2369] = 8'h00;
    mem[2370] = 8'h00;
    mem[2371] = 8'h00;
    mem[2372] = 8'hfc;
    mem[2373] = 8'h01;
    mem[2374] = 8'hf8;
    mem[2375] = 8'h1f;
    mem[2376] = 8'h00;
    mem[2377] = 8'hf0;
    mem[2378] = 8'h03;
    mem[2379] = 8'hf8;
    mem[2380] = 8'h7f;
    mem[2381] = 8'h00;
    mem[2382] = 8'h00;
    mem[2383] = 8'h70;
    mem[2384] = 8'h00;
    mem[2385] = 8'h00;
    mem[2386] = 8'hc0;
    mem[2387] = 8'hdf;
    mem[2388] = 8'hff;
    mem[2389] = 8'h3f;
    mem[2390] = 8'h00;
    mem[2391] = 8'hc0;
    mem[2392] = 8'hff;
    mem[2393] = 8'h01;
    mem[2394] = 8'hfc;
    mem[2395] = 8'h03;
    mem[2396] = 8'h00;
    mem[2397] = 8'h00;
    mem[2398] = 8'h00;
    mem[2399] = 8'h00;
    mem[2400] = 8'h00;
    mem[2401] = 8'h00;
    mem[2402] = 8'h00;
    mem[2403] = 8'h00;
    mem[2404] = 8'hfe;
    mem[2405] = 8'h01;
    mem[2406] = 8'hfc;
    mem[2407] = 8'h0f;
    mem[2408] = 8'h00;
    mem[2409] = 8'hf8;
    mem[2410] = 8'h00;
    mem[2411] = 8'hf0;
    mem[2412] = 8'h3f;
    mem[2413] = 8'h00;
    mem[2414] = 8'h00;
    mem[2415] = 8'h70;
    mem[2416] = 8'h00;
    mem[2417] = 8'h00;
    mem[2418] = 8'h00;
    mem[2419] = 8'h80;
    mem[2420] = 8'hff;
    mem[2421] = 8'h7f;
    mem[2422] = 8'h00;
    mem[2423] = 8'h00;
    mem[2424] = 8'hff;
    mem[2425] = 8'h01;
    mem[2426] = 8'hfc;
    mem[2427] = 8'h03;
    mem[2428] = 8'h00;
    mem[2429] = 8'h00;
    mem[2430] = 8'h00;
    mem[2431] = 8'h00;
    mem[2432] = 8'h00;
    mem[2433] = 8'h00;
    mem[2434] = 8'h00;
    mem[2435] = 8'h00;
    mem[2436] = 8'hfe;
    mem[2437] = 8'h01;
    mem[2438] = 8'hfc;
    mem[2439] = 8'h03;
    mem[2440] = 8'h00;
    mem[2441] = 8'h7e;
    mem[2442] = 8'h00;
    mem[2443] = 8'hf8;
    mem[2444] = 8'h1f;
    mem[2445] = 8'h00;
    mem[2446] = 8'h00;
    mem[2447] = 8'h70;
    mem[2448] = 8'h00;
    mem[2449] = 8'h00;
    mem[2450] = 8'h00;
    mem[2451] = 8'h00;
    mem[2452] = 8'hfe;
    mem[2453] = 8'hff;
    mem[2454] = 8'h01;
    mem[2455] = 8'h00;
    mem[2456] = 8'hfe;
    mem[2457] = 8'h01;
    mem[2458] = 8'hfc;
    mem[2459] = 8'h03;
    mem[2460] = 8'h00;
    mem[2461] = 8'h00;
    mem[2462] = 8'h00;
    mem[2463] = 8'h00;
    mem[2464] = 8'h00;
    mem[2465] = 8'h00;
    mem[2466] = 8'h00;
    mem[2467] = 8'h00;
    mem[2468] = 8'hfe;
    mem[2469] = 8'h01;
    mem[2470] = 8'hfc;
    mem[2471] = 8'h03;
    mem[2472] = 8'he0;
    mem[2473] = 8'h1f;
    mem[2474] = 8'h00;
    mem[2475] = 8'h7e;
    mem[2476] = 8'h00;
    mem[2477] = 8'h00;
    mem[2478] = 8'h00;
    mem[2479] = 8'h70;
    mem[2480] = 8'h00;
    mem[2481] = 8'h00;
    mem[2482] = 8'h00;
    mem[2483] = 8'h00;
    mem[2484] = 8'hf8;
    mem[2485] = 8'hff;
    mem[2486] = 8'h03;
    mem[2487] = 8'h00;
    mem[2488] = 8'hfc;
    mem[2489] = 8'h01;
    mem[2490] = 8'hf8;
    mem[2491] = 8'h03;
    mem[2492] = 8'h00;
    mem[2493] = 8'h00;
    mem[2494] = 8'h00;
    mem[2495] = 8'h00;
    mem[2496] = 8'h00;
    mem[2497] = 8'h00;
    mem[2498] = 8'h00;
    mem[2499] = 8'h00;
    mem[2500] = 8'hfe;
    mem[2501] = 8'h01;
    mem[2502] = 8'hfc;
    mem[2503] = 8'h03;
    mem[2504] = 8'hf8;
    mem[2505] = 8'h0f;
    mem[2506] = 8'h00;
    mem[2507] = 8'h1f;
    mem[2508] = 8'h00;
    mem[2509] = 8'h00;
    mem[2510] = 8'h00;
    mem[2511] = 8'h70;
    mem[2512] = 8'h00;
    mem[2513] = 8'h00;
    mem[2514] = 8'h00;
    mem[2515] = 8'h00;
    mem[2516] = 8'hf0;
    mem[2517] = 8'hff;
    mem[2518] = 8'h0f;
    mem[2519] = 8'h00;
    mem[2520] = 8'hfc;
    mem[2521] = 8'h03;
    mem[2522] = 8'hf8;
    mem[2523] = 8'h03;
    mem[2524] = 8'h00;
    mem[2525] = 8'h00;
    mem[2526] = 8'h00;
    mem[2527] = 8'h00;
    mem[2528] = 8'h00;
    mem[2529] = 8'h00;
    mem[2530] = 8'h00;
    mem[2531] = 8'h00;
    mem[2532] = 8'hfe;
    mem[2533] = 8'h01;
    mem[2534] = 8'hfc;
    mem[2535] = 8'h01;
    mem[2536] = 8'hfe;
    mem[2537] = 8'h1f;
    mem[2538] = 8'hc0;
    mem[2539] = 8'h0f;
    mem[2540] = 8'h00;
    mem[2541] = 8'h00;
    mem[2542] = 8'h00;
    mem[2543] = 8'h00;
    mem[2544] = 8'h00;
    mem[2545] = 8'h00;
    mem[2546] = 8'h00;
    mem[2547] = 8'h00;
    mem[2548] = 8'hc0;
    mem[2549] = 8'hff;
    mem[2550] = 8'h1f;
    mem[2551] = 8'h00;
    mem[2552] = 8'hfc;
    mem[2553] = 8'h03;
    mem[2554] = 8'hf8;
    mem[2555] = 8'h03;
    mem[2556] = 8'h00;
    mem[2557] = 8'h00;
    mem[2558] = 8'h00;
    mem[2559] = 8'h00;
    mem[2560] = 8'h00;
    mem[2561] = 8'h00;
    mem[2562] = 8'h00;
    mem[2563] = 8'h00;
    mem[2564] = 8'hfe;
    mem[2565] = 8'h01;
    mem[2566] = 8'hfc;
    mem[2567] = 8'h01;
    mem[2568] = 8'h3e;
    mem[2569] = 8'h3e;
    mem[2570] = 8'he0;
    mem[2571] = 8'h03;
    mem[2572] = 8'h00;
    mem[2573] = 8'h00;
    mem[2574] = 8'h00;
    mem[2575] = 8'h00;
    mem[2576] = 8'h00;
    mem[2577] = 8'h00;
    mem[2578] = 8'h00;
    mem[2579] = 8'h00;
    mem[2580] = 8'h00;
    mem[2581] = 8'hff;
    mem[2582] = 8'h7f;
    mem[2583] = 8'h00;
    mem[2584] = 8'hfc;
    mem[2585] = 8'h03;
    mem[2586] = 8'hf8;
    mem[2587] = 8'h03;
    mem[2588] = 8'h00;
    mem[2589] = 8'h00;
    mem[2590] = 8'h00;
    mem[2591] = 8'h00;
    mem[2592] = 8'h00;
    mem[2593] = 8'h00;
    mem[2594] = 8'h00;
    mem[2595] = 8'h00;
    mem[2596] = 8'hfe;
    mem[2597] = 8'h01;
    mem[2598] = 8'hfc;
    mem[2599] = 8'h01;
    mem[2600] = 8'h0f;
    mem[2601] = 8'h78;
    mem[2602] = 8'hf8;
    mem[2603] = 8'h01;
    mem[2604] = 8'h00;
    mem[2605] = 8'h00;
    mem[2606] = 8'h00;
    mem[2607] = 8'h00;
    mem[2608] = 8'h00;
    mem[2609] = 8'h00;
    mem[2610] = 8'h00;
    mem[2611] = 8'h00;
    mem[2612] = 8'h00;
    mem[2613] = 8'hfe;
    mem[2614] = 8'hff;
    mem[2615] = 8'h00;
    mem[2616] = 8'hfc;
    mem[2617] = 8'h03;
    mem[2618] = 8'hf8;
    mem[2619] = 8'h03;
    mem[2620] = 8'h00;
    mem[2621] = 8'h00;
    mem[2622] = 8'h00;
    mem[2623] = 8'h00;
    mem[2624] = 8'h00;
    mem[2625] = 8'h00;
    mem[2626] = 8'h00;
    mem[2627] = 8'h00;
    mem[2628] = 8'hfe;
    mem[2629] = 8'h01;
    mem[2630] = 8'hfc;
    mem[2631] = 8'h01;
    mem[2632] = 8'he7;
    mem[2633] = 8'h73;
    mem[2634] = 8'h7c;
    mem[2635] = 8'h00;
    mem[2636] = 8'h00;
    mem[2637] = 8'hf0;
    mem[2638] = 8'hff;
    mem[2639] = 8'hff;
    mem[2640] = 8'hff;
    mem[2641] = 8'h03;
    mem[2642] = 8'h00;
    mem[2643] = 8'h00;
    mem[2644] = 8'h00;
    mem[2645] = 8'hf8;
    mem[2646] = 8'hff;
    mem[2647] = 8'h01;
    mem[2648] = 8'hfc;
    mem[2649] = 8'h03;
    mem[2650] = 8'hf8;
    mem[2651] = 8'h03;
    mem[2652] = 8'h00;
    mem[2653] = 8'h00;
    mem[2654] = 8'h00;
    mem[2655] = 8'h00;
    mem[2656] = 8'h00;
    mem[2657] = 8'h00;
    mem[2658] = 8'h00;
    mem[2659] = 8'h00;
    mem[2660] = 8'hfe;
    mem[2661] = 8'h01;
    mem[2662] = 8'hfc;
    mem[2663] = 8'h81;
    mem[2664] = 8'hf3;
    mem[2665] = 8'hf7;
    mem[2666] = 8'h3f;
    mem[2667] = 8'h00;
    mem[2668] = 8'h00;
    mem[2669] = 8'hf8;
    mem[2670] = 8'hff;
    mem[2671] = 8'hff;
    mem[2672] = 8'hff;
    mem[2673] = 8'h3f;
    mem[2674] = 8'h00;
    mem[2675] = 8'h00;
    mem[2676] = 8'h00;
    mem[2677] = 8'he0;
    mem[2678] = 8'hff;
    mem[2679] = 8'h01;
    mem[2680] = 8'hf8;
    mem[2681] = 8'h03;
    mem[2682] = 8'hf8;
    mem[2683] = 8'h07;
    mem[2684] = 8'h00;
    mem[2685] = 8'h00;
    mem[2686] = 8'h00;
    mem[2687] = 8'h00;
    mem[2688] = 8'h00;
    mem[2689] = 8'h00;
    mem[2690] = 8'h00;
    mem[2691] = 8'h00;
    mem[2692] = 8'hfe;
    mem[2693] = 8'h01;
    mem[2694] = 8'hfe;
    mem[2695] = 8'h81;
    mem[2696] = 8'hf3;
    mem[2697] = 8'he7;
    mem[2698] = 8'h0f;
    mem[2699] = 8'h00;
    mem[2700] = 8'h00;
    mem[2701] = 8'hfc;
    mem[2702] = 8'hff;
    mem[2703] = 8'hff;
    mem[2704] = 8'hff;
    mem[2705] = 8'hff;
    mem[2706] = 8'h00;
    mem[2707] = 8'h00;
    mem[2708] = 8'h00;
    mem[2709] = 8'he0;
    mem[2710] = 8'hff;
    mem[2711] = 8'h03;
    mem[2712] = 8'hf8;
    mem[2713] = 8'h03;
    mem[2714] = 8'hf8;
    mem[2715] = 8'h07;
    mem[2716] = 8'h00;
    mem[2717] = 8'h00;
    mem[2718] = 8'h00;
    mem[2719] = 8'h00;
    mem[2720] = 8'h00;
    mem[2721] = 8'h00;
    mem[2722] = 8'h00;
    mem[2723] = 8'h00;
    mem[2724] = 8'hfe;
    mem[2725] = 8'h01;
    mem[2726] = 8'hfe;
    mem[2727] = 8'h81;
    mem[2728] = 8'h3b;
    mem[2729] = 8'he7;
    mem[2730] = 8'h07;
    mem[2731] = 8'h00;
    mem[2732] = 8'h00;
    mem[2733] = 8'hfe;
    mem[2734] = 8'hff;
    mem[2735] = 8'hff;
    mem[2736] = 8'hff;
    mem[2737] = 8'hff;
    mem[2738] = 8'h03;
    mem[2739] = 8'h00;
    mem[2740] = 8'h00;
    mem[2741] = 8'he0;
    mem[2742] = 8'hff;
    mem[2743] = 8'h03;
    mem[2744] = 8'hf8;
    mem[2745] = 8'h03;
    mem[2746] = 8'hf8;
    mem[2747] = 8'h07;
    mem[2748] = 8'h00;
    mem[2749] = 8'h00;
    mem[2750] = 8'h00;
    mem[2751] = 8'h00;
    mem[2752] = 8'h00;
    mem[2753] = 8'h00;
    mem[2754] = 8'h00;
    mem[2755] = 8'h00;
    mem[2756] = 8'hfe;
    mem[2757] = 8'h01;
    mem[2758] = 8'hfe;
    mem[2759] = 8'h81;
    mem[2760] = 8'h7b;
    mem[2761] = 8'he7;
    mem[2762] = 8'h01;
    mem[2763] = 8'h00;
    mem[2764] = 8'h00;
    mem[2765] = 8'hfe;
    mem[2766] = 8'hff;
    mem[2767] = 8'hff;
    mem[2768] = 8'hff;
    mem[2769] = 8'hff;
    mem[2770] = 8'h07;
    mem[2771] = 8'h00;
    mem[2772] = 8'h00;
    mem[2773] = 8'he0;
    mem[2774] = 8'hfe;
    mem[2775] = 8'h07;
    mem[2776] = 8'hf8;
    mem[2777] = 8'h03;
    mem[2778] = 8'hf8;
    mem[2779] = 8'h07;
    mem[2780] = 8'h00;
    mem[2781] = 8'h00;
    mem[2782] = 8'h00;
    mem[2783] = 8'h00;
    mem[2784] = 8'h00;
    mem[2785] = 8'h00;
    mem[2786] = 8'h00;
    mem[2787] = 8'h00;
    mem[2788] = 8'hfe;
    mem[2789] = 8'h00;
    mem[2790] = 8'hfe;
    mem[2791] = 8'h81;
    mem[2792] = 8'hf3;
    mem[2793] = 8'hf7;
    mem[2794] = 8'h00;
    mem[2795] = 8'h00;
    mem[2796] = 8'h00;
    mem[2797] = 8'hfe;
    mem[2798] = 8'hff;
    mem[2799] = 8'hff;
    mem[2800] = 8'hff;
    mem[2801] = 8'hff;
    mem[2802] = 8'h0f;
    mem[2803] = 8'h00;
    mem[2804] = 8'h00;
    mem[2805] = 8'he0;
    mem[2806] = 8'hf8;
    mem[2807] = 8'h07;
    mem[2808] = 8'hf8;
    mem[2809] = 8'h03;
    mem[2810] = 8'hf8;
    mem[2811] = 8'h07;
    mem[2812] = 8'h00;
    mem[2813] = 8'h00;
    mem[2814] = 8'h00;
    mem[2815] = 8'h00;
    mem[2816] = 8'h00;
    mem[2817] = 8'h00;
    mem[2818] = 8'h00;
    mem[2819] = 8'h00;
    mem[2820] = 8'hfe;
    mem[2821] = 8'h00;
    mem[2822] = 8'hfe;
    mem[2823] = 8'h81;
    mem[2824] = 8'he7;
    mem[2825] = 8'h73;
    mem[2826] = 8'h00;
    mem[2827] = 8'h00;
    mem[2828] = 8'h00;
    mem[2829] = 8'hfe;
    mem[2830] = 8'hff;
    mem[2831] = 8'hff;
    mem[2832] = 8'hff;
    mem[2833] = 8'hff;
    mem[2834] = 8'h0f;
    mem[2835] = 8'h00;
    mem[2836] = 8'h00;
    mem[2837] = 8'he0;
    mem[2838] = 8'he0;
    mem[2839] = 8'h07;
    mem[2840] = 8'hf8;
    mem[2841] = 8'h03;
    mem[2842] = 8'hf8;
    mem[2843] = 8'h07;
    mem[2844] = 8'h00;
    mem[2845] = 8'h00;
    mem[2846] = 8'h00;
    mem[2847] = 8'h00;
    mem[2848] = 8'h00;
    mem[2849] = 8'h00;
    mem[2850] = 8'h00;
    mem[2851] = 8'h00;
    mem[2852] = 8'hfe;
    mem[2853] = 8'h00;
    mem[2854] = 8'hfe;
    mem[2855] = 8'h01;
    mem[2856] = 8'hcf;
    mem[2857] = 8'h79;
    mem[2858] = 8'h00;
    mem[2859] = 8'h00;
    mem[2860] = 8'h00;
    mem[2861] = 8'hfe;
    mem[2862] = 8'hff;
    mem[2863] = 8'hff;
    mem[2864] = 8'hff;
    mem[2865] = 8'hff;
    mem[2866] = 8'h1f;
    mem[2867] = 8'h00;
    mem[2868] = 8'h00;
    mem[2869] = 8'he0;
    mem[2870] = 8'hc0;
    mem[2871] = 8'h07;
    mem[2872] = 8'hf8;
    mem[2873] = 8'h03;
    mem[2874] = 8'hf8;
    mem[2875] = 8'h07;
    mem[2876] = 8'h00;
    mem[2877] = 8'h00;
    mem[2878] = 8'h00;
    mem[2879] = 8'h00;
    mem[2880] = 8'h00;
    mem[2881] = 8'h00;
    mem[2882] = 8'h00;
    mem[2883] = 8'h00;
    mem[2884] = 8'hfe;
    mem[2885] = 8'h00;
    mem[2886] = 8'hfe;
    mem[2887] = 8'h01;
    mem[2888] = 8'h1f;
    mem[2889] = 8'h7c;
    mem[2890] = 8'h00;
    mem[2891] = 8'h00;
    mem[2892] = 8'h00;
    mem[2893] = 8'hfe;
    mem[2894] = 8'hff;
    mem[2895] = 8'hff;
    mem[2896] = 8'hff;
    mem[2897] = 8'hff;
    mem[2898] = 8'h3f;
    mem[2899] = 8'h00;
    mem[2900] = 8'h00;
    mem[2901] = 8'he0;
    mem[2902] = 8'h00;
    mem[2903] = 8'h07;
    mem[2904] = 8'hf8;
    mem[2905] = 8'h03;
    mem[2906] = 8'hfe;
    mem[2907] = 8'h0f;
    mem[2908] = 8'h00;
    mem[2909] = 8'h00;
    mem[2910] = 8'h00;
    mem[2911] = 8'h00;
    mem[2912] = 8'h00;
    mem[2913] = 8'h00;
    mem[2914] = 8'h00;
    mem[2915] = 8'h00;
    mem[2916] = 8'hfe;
    mem[2917] = 8'h00;
    mem[2918] = 8'hfe;
    mem[2919] = 8'h01;
    mem[2920] = 8'hff;
    mem[2921] = 8'h7f;
    mem[2922] = 8'h00;
    mem[2923] = 8'h00;
    mem[2924] = 8'h00;
    mem[2925] = 8'hfe;
    mem[2926] = 8'hff;
    mem[2927] = 8'hff;
    mem[2928] = 8'hff;
    mem[2929] = 8'hff;
    mem[2930] = 8'h3f;
    mem[2931] = 8'h00;
    mem[2932] = 8'h00;
    mem[2933] = 8'he0;
    mem[2934] = 8'h00;
    mem[2935] = 8'h07;
    mem[2936] = 8'hf8;
    mem[2937] = 8'h07;
    mem[2938] = 8'hfe;
    mem[2939] = 8'h1f;
    mem[2940] = 8'h00;
    mem[2941] = 8'h00;
    mem[2942] = 8'h00;
    mem[2943] = 8'h00;
    mem[2944] = 8'h00;
    mem[2945] = 8'h00;
    mem[2946] = 8'h00;
    mem[2947] = 8'h00;
    mem[2948] = 8'hfe;
    mem[2949] = 8'h00;
    mem[2950] = 8'hfe;
    mem[2951] = 8'h01;
    mem[2952] = 8'hff;
    mem[2953] = 8'h7f;
    mem[2954] = 8'h00;
    mem[2955] = 8'h00;
    mem[2956] = 8'h00;
    mem[2957] = 8'hfe;
    mem[2958] = 8'h1f;
    mem[2959] = 8'h00;
    mem[2960] = 8'h80;
    mem[2961] = 8'hff;
    mem[2962] = 8'h3f;
    mem[2963] = 8'h00;
    mem[2964] = 8'h00;
    mem[2965] = 8'he0;
    mem[2966] = 8'h00;
    mem[2967] = 8'h07;
    mem[2968] = 8'hf8;
    mem[2969] = 8'h07;
    mem[2970] = 8'hff;
    mem[2971] = 8'h3f;
    mem[2972] = 8'h00;
    mem[2973] = 8'h00;
    mem[2974] = 8'h00;
    mem[2975] = 8'h00;
    mem[2976] = 8'h00;
    mem[2977] = 8'h00;
    mem[2978] = 8'h00;
    mem[2979] = 8'h00;
    mem[2980] = 8'hfe;
    mem[2981] = 8'h00;
    mem[2982] = 8'hfe;
    mem[2983] = 8'h01;
    mem[2984] = 8'hff;
    mem[2985] = 8'h77;
    mem[2986] = 8'h00;
    mem[2987] = 8'h00;
    mem[2988] = 8'h00;
    mem[2989] = 8'hfe;
    mem[2990] = 8'h1f;
    mem[2991] = 8'h00;
    mem[2992] = 8'h00;
    mem[2993] = 8'hfe;
    mem[2994] = 8'h7f;
    mem[2995] = 8'h00;
    mem[2996] = 8'h00;
    mem[2997] = 8'he0;
    mem[2998] = 8'h00;
    mem[2999] = 8'h07;
    mem[3000] = 8'hf8;
    mem[3001] = 8'h87;
    mem[3002] = 8'h3f;
    mem[3003] = 8'h7f;
    mem[3004] = 8'h00;
    mem[3005] = 8'h00;
    mem[3006] = 8'h00;
    mem[3007] = 8'h00;
    mem[3008] = 8'h00;
    mem[3009] = 8'h00;
    mem[3010] = 8'h00;
    mem[3011] = 8'h00;
    mem[3012] = 8'hfe;
    mem[3013] = 8'h00;
    mem[3014] = 8'hfe;
    mem[3015] = 8'h01;
    mem[3016] = 8'h0f;
    mem[3017] = 8'h70;
    mem[3018] = 8'h00;
    mem[3019] = 8'h00;
    mem[3020] = 8'h00;
    mem[3021] = 8'hfe;
    mem[3022] = 8'h1f;
    mem[3023] = 8'h00;
    mem[3024] = 8'h00;
    mem[3025] = 8'hfc;
    mem[3026] = 8'h7f;
    mem[3027] = 8'h00;
    mem[3028] = 8'h00;
    mem[3029] = 8'he0;
    mem[3030] = 8'h00;
    mem[3031] = 8'h07;
    mem[3032] = 8'hf8;
    mem[3033] = 8'h87;
    mem[3034] = 8'h0f;
    mem[3035] = 8'h7c;
    mem[3036] = 8'h00;
    mem[3037] = 8'h00;
    mem[3038] = 8'h00;
    mem[3039] = 8'h00;
    mem[3040] = 8'h00;
    mem[3041] = 8'h00;
    mem[3042] = 8'h00;
    mem[3043] = 8'h00;
    mem[3044] = 8'hfe;
    mem[3045] = 8'h00;
    mem[3046] = 8'hfe;
    mem[3047] = 8'h01;
    mem[3048] = 8'h0f;
    mem[3049] = 8'h70;
    mem[3050] = 8'h00;
    mem[3051] = 8'h00;
    mem[3052] = 8'h00;
    mem[3053] = 8'hfe;
    mem[3054] = 8'h1f;
    mem[3055] = 8'h00;
    mem[3056] = 8'h00;
    mem[3057] = 8'hfc;
    mem[3058] = 8'h7f;
    mem[3059] = 8'h00;
    mem[3060] = 8'h00;
    mem[3061] = 8'he0;
    mem[3062] = 8'h00;
    mem[3063] = 8'h07;
    mem[3064] = 8'hf8;
    mem[3065] = 8'hc7;
    mem[3066] = 8'h07;
    mem[3067] = 8'hf8;
    mem[3068] = 8'h00;
    mem[3069] = 8'h00;
    mem[3070] = 8'h00;
    mem[3071] = 8'h00;
    mem[3072] = 8'h00;
    mem[3073] = 8'h00;
    mem[3074] = 8'h00;
    mem[3075] = 8'h00;
    mem[3076] = 8'hfe;
    mem[3077] = 8'h00;
    mem[3078] = 8'hfe;
    mem[3079] = 8'h01;
    mem[3080] = 8'h0f;
    mem[3081] = 8'h70;
    mem[3082] = 8'h00;
    mem[3083] = 8'h00;
    mem[3084] = 8'h00;
    mem[3085] = 8'hfe;
    mem[3086] = 8'h1f;
    mem[3087] = 8'h00;
    mem[3088] = 8'h00;
    mem[3089] = 8'hf8;
    mem[3090] = 8'h7f;
    mem[3091] = 8'h00;
    mem[3092] = 8'h00;
    mem[3093] = 8'he0;
    mem[3094] = 8'h00;
    mem[3095] = 8'h07;
    mem[3096] = 8'hf8;
    mem[3097] = 8'hc7;
    mem[3098] = 8'h07;
    mem[3099] = 8'hf8;
    mem[3100] = 8'h00;
    mem[3101] = 8'h00;
    mem[3102] = 8'h00;
    mem[3103] = 8'h00;
    mem[3104] = 8'h00;
    mem[3105] = 8'h00;
    mem[3106] = 8'h00;
    mem[3107] = 8'h00;
    mem[3108] = 8'hff;
    mem[3109] = 8'h00;
    mem[3110] = 8'hfe;
    mem[3111] = 8'h00;
    mem[3112] = 8'h0f;
    mem[3113] = 8'h70;
    mem[3114] = 8'h00;
    mem[3115] = 8'h00;
    mem[3116] = 8'h00;
    mem[3117] = 8'hfe;
    mem[3118] = 8'h1f;
    mem[3119] = 8'h00;
    mem[3120] = 8'h00;
    mem[3121] = 8'hf8;
    mem[3122] = 8'h7f;
    mem[3123] = 8'h00;
    mem[3124] = 8'h00;
    mem[3125] = 8'he0;
    mem[3126] = 8'h00;
    mem[3127] = 8'h07;
    mem[3128] = 8'hf8;
    mem[3129] = 8'hc7;
    mem[3130] = 8'h07;
    mem[3131] = 8'hf8;
    mem[3132] = 8'h00;
    mem[3133] = 8'h00;
    mem[3134] = 8'h00;
    mem[3135] = 8'h00;
    mem[3136] = 8'h00;
    mem[3137] = 8'h00;
    mem[3138] = 8'h00;
    mem[3139] = 8'h00;
    mem[3140] = 8'hff;
    mem[3141] = 8'h00;
    mem[3142] = 8'hfe;
    mem[3143] = 8'h00;
    mem[3144] = 8'h0f;
    mem[3145] = 8'h70;
    mem[3146] = 8'h00;
    mem[3147] = 8'h00;
    mem[3148] = 8'h00;
    mem[3149] = 8'hfe;
    mem[3150] = 8'h1f;
    mem[3151] = 8'h00;
    mem[3152] = 8'h00;
    mem[3153] = 8'hf8;
    mem[3154] = 8'h7f;
    mem[3155] = 8'h00;
    mem[3156] = 8'h00;
    mem[3157] = 8'he0;
    mem[3158] = 8'h00;
    mem[3159] = 8'h07;
    mem[3160] = 8'hf8;
    mem[3161] = 8'hc7;
    mem[3162] = 8'h07;
    mem[3163] = 8'hf8;
    mem[3164] = 8'h00;
    mem[3165] = 8'h00;
    mem[3166] = 8'h00;
    mem[3167] = 8'h00;
    mem[3168] = 8'h00;
    mem[3169] = 8'h00;
    mem[3170] = 8'h00;
    mem[3171] = 8'h00;
    mem[3172] = 8'hff;
    mem[3173] = 8'h00;
    mem[3174] = 8'hfe;
    mem[3175] = 8'h00;
    mem[3176] = 8'h0f;
    mem[3177] = 8'h70;
    mem[3178] = 8'h00;
    mem[3179] = 8'h00;
    mem[3180] = 8'h00;
    mem[3181] = 8'hfe;
    mem[3182] = 8'h1f;
    mem[3183] = 8'h00;
    mem[3184] = 8'h00;
    mem[3185] = 8'hf8;
    mem[3186] = 8'h7f;
    mem[3187] = 8'h00;
    mem[3188] = 8'h00;
    mem[3189] = 8'he0;
    mem[3190] = 8'h00;
    mem[3191] = 8'h07;
    mem[3192] = 8'hf8;
    mem[3193] = 8'h87;
    mem[3194] = 8'h0f;
    mem[3195] = 8'h7c;
    mem[3196] = 8'h00;
    mem[3197] = 8'h00;
    mem[3198] = 8'h00;
    mem[3199] = 8'h00;
    mem[3200] = 8'h00;
    mem[3201] = 8'h00;
    mem[3202] = 8'h00;
    mem[3203] = 8'h00;
    mem[3204] = 8'hff;
    mem[3205] = 8'h00;
    mem[3206] = 8'hfe;
    mem[3207] = 8'h00;
    mem[3208] = 8'h0f;
    mem[3209] = 8'h70;
    mem[3210] = 8'h00;
    mem[3211] = 8'h00;
    mem[3212] = 8'h00;
    mem[3213] = 8'hfe;
    mem[3214] = 8'h1f;
    mem[3215] = 8'h00;
    mem[3216] = 8'h00;
    mem[3217] = 8'hf8;
    mem[3218] = 8'h7f;
    mem[3219] = 8'h00;
    mem[3220] = 8'h00;
    mem[3221] = 8'he0;
    mem[3222] = 8'h00;
    mem[3223] = 8'h07;
    mem[3224] = 8'hf8;
    mem[3225] = 8'h87;
    mem[3226] = 8'h0f;
    mem[3227] = 8'h7e;
    mem[3228] = 8'h00;
    mem[3229] = 8'h00;
    mem[3230] = 8'h00;
    mem[3231] = 8'h00;
    mem[3232] = 8'h00;
    mem[3233] = 8'h00;
    mem[3234] = 8'h00;
    mem[3235] = 8'h00;
    mem[3236] = 8'hff;
    mem[3237] = 8'h00;
    mem[3238] = 8'hfe;
    mem[3239] = 8'h00;
    mem[3240] = 8'h0f;
    mem[3241] = 8'h70;
    mem[3242] = 8'h00;
    mem[3243] = 8'h00;
    mem[3244] = 8'h00;
    mem[3245] = 8'hfe;
    mem[3246] = 8'h1f;
    mem[3247] = 8'h00;
    mem[3248] = 8'h00;
    mem[3249] = 8'hf8;
    mem[3250] = 8'h7f;
    mem[3251] = 8'h00;
    mem[3252] = 8'h00;
    mem[3253] = 8'he0;
    mem[3254] = 8'h00;
    mem[3255] = 8'h07;
    mem[3256] = 8'hf8;
    mem[3257] = 8'h87;
    mem[3258] = 8'hff;
    mem[3259] = 8'h7f;
    mem[3260] = 8'h00;
    mem[3261] = 8'h00;
    mem[3262] = 8'h00;
    mem[3263] = 8'h00;
    mem[3264] = 8'h00;
    mem[3265] = 8'h00;
    mem[3266] = 8'h00;
    mem[3267] = 8'h00;
    mem[3268] = 8'hff;
    mem[3269] = 8'h00;
    mem[3270] = 8'hfe;
    mem[3271] = 8'h00;
    mem[3272] = 8'h0f;
    mem[3273] = 8'h70;
    mem[3274] = 8'h00;
    mem[3275] = 8'h00;
    mem[3276] = 8'h00;
    mem[3277] = 8'hfe;
    mem[3278] = 8'h1f;
    mem[3279] = 8'h00;
    mem[3280] = 8'h00;
    mem[3281] = 8'hf8;
    mem[3282] = 8'h7f;
    mem[3283] = 8'h00;
    mem[3284] = 8'h00;
    mem[3285] = 8'he0;
    mem[3286] = 8'h00;
    mem[3287] = 8'h07;
    mem[3288] = 8'hf8;
    mem[3289] = 8'h07;
    mem[3290] = 8'hff;
    mem[3291] = 8'h3f;
    mem[3292] = 8'h00;
    mem[3293] = 8'h00;
    mem[3294] = 8'h00;
    mem[3295] = 8'h00;
    mem[3296] = 8'h00;
    mem[3297] = 8'h00;
    mem[3298] = 8'h00;
    mem[3299] = 8'h00;
    mem[3300] = 8'hff;
    mem[3301] = 8'h00;
    mem[3302] = 8'hfe;
    mem[3303] = 8'h00;
    mem[3304] = 8'h0f;
    mem[3305] = 8'h70;
    mem[3306] = 8'h00;
    mem[3307] = 8'h00;
    mem[3308] = 8'h00;
    mem[3309] = 8'hfe;
    mem[3310] = 8'h1f;
    mem[3311] = 8'h00;
    mem[3312] = 8'h00;
    mem[3313] = 8'hf8;
    mem[3314] = 8'h3f;
    mem[3315] = 8'h00;
    mem[3316] = 8'h00;
    mem[3317] = 8'he0;
    mem[3318] = 8'h00;
    mem[3319] = 8'h07;
    mem[3320] = 8'hf8;
    mem[3321] = 8'h07;
    mem[3322] = 8'hfe;
    mem[3323] = 8'h1f;
    mem[3324] = 8'h00;
    mem[3325] = 8'h00;
    mem[3326] = 8'h00;
    mem[3327] = 8'h00;
    mem[3328] = 8'h00;
    mem[3329] = 8'h00;
    mem[3330] = 8'h00;
    mem[3331] = 8'h00;
    mem[3332] = 8'hff;
    mem[3333] = 8'h00;
    mem[3334] = 8'hfe;
    mem[3335] = 8'h00;
    mem[3336] = 8'h0f;
    mem[3337] = 8'h70;
    mem[3338] = 8'h00;
    mem[3339] = 8'h00;
    mem[3340] = 8'h00;
    mem[3341] = 8'hfe;
    mem[3342] = 8'h1f;
    mem[3343] = 8'h00;
    mem[3344] = 8'h00;
    mem[3345] = 8'hfc;
    mem[3346] = 8'h3f;
    mem[3347] = 8'h00;
    mem[3348] = 8'h00;
    mem[3349] = 8'he0;
    mem[3350] = 8'h00;
    mem[3351] = 8'h07;
    mem[3352] = 8'hf8;
    mem[3353] = 8'h07;
    mem[3354] = 8'hfc;
    mem[3355] = 8'h0f;
    mem[3356] = 8'h00;
    mem[3357] = 8'h00;
    mem[3358] = 8'h00;
    mem[3359] = 8'h00;
    mem[3360] = 8'h00;
    mem[3361] = 8'h00;
    mem[3362] = 8'h00;
    mem[3363] = 8'h00;
    mem[3364] = 8'hff;
    mem[3365] = 8'h00;
    mem[3366] = 8'hfe;
    mem[3367] = 8'h00;
    mem[3368] = 8'h0f;
    mem[3369] = 8'h70;
    mem[3370] = 8'h00;
    mem[3371] = 8'h00;
    mem[3372] = 8'h00;
    mem[3373] = 8'hfe;
    mem[3374] = 8'h1f;
    mem[3375] = 8'h00;
    mem[3376] = 8'h00;
    mem[3377] = 8'hfe;
    mem[3378] = 8'h3f;
    mem[3379] = 8'h00;
    mem[3380] = 8'h00;
    mem[3381] = 8'he0;
    mem[3382] = 8'h00;
    mem[3383] = 8'h07;
    mem[3384] = 8'hf8;
    mem[3385] = 8'h07;
    mem[3386] = 8'hf0;
    mem[3387] = 8'h03;
    mem[3388] = 8'h00;
    mem[3389] = 8'h00;
    mem[3390] = 8'h00;
    mem[3391] = 8'h00;
    mem[3392] = 8'h00;
    mem[3393] = 8'h00;
    mem[3394] = 8'h00;
    mem[3395] = 8'h00;
    mem[3396] = 8'hff;
    mem[3397] = 8'h00;
    mem[3398] = 8'hfe;
    mem[3399] = 8'h00;
    mem[3400] = 8'h0f;
    mem[3401] = 8'h70;
    mem[3402] = 8'h00;
    mem[3403] = 8'h00;
    mem[3404] = 8'h00;
    mem[3405] = 8'hfe;
    mem[3406] = 8'h1f;
    mem[3407] = 8'h00;
    mem[3408] = 8'h80;
    mem[3409] = 8'hff;
    mem[3410] = 8'h1f;
    mem[3411] = 8'h00;
    mem[3412] = 8'h00;
    mem[3413] = 8'he0;
    mem[3414] = 8'h00;
    mem[3415] = 8'h07;
    mem[3416] = 8'hf8;
    mem[3417] = 8'h07;
    mem[3418] = 8'h00;
    mem[3419] = 8'h00;
    mem[3420] = 8'h00;
    mem[3421] = 8'h00;
    mem[3422] = 8'h00;
    mem[3423] = 8'h00;
    mem[3424] = 8'h00;
    mem[3425] = 8'h00;
    mem[3426] = 8'h00;
    mem[3427] = 8'h00;
    mem[3428] = 8'hff;
    mem[3429] = 8'h00;
    mem[3430] = 8'hfe;
    mem[3431] = 8'h00;
    mem[3432] = 8'h0f;
    mem[3433] = 8'h70;
    mem[3434] = 8'h00;
    mem[3435] = 8'h00;
    mem[3436] = 8'h00;
    mem[3437] = 8'hfe;
    mem[3438] = 8'hff;
    mem[3439] = 8'hff;
    mem[3440] = 8'hff;
    mem[3441] = 8'hff;
    mem[3442] = 8'h1f;
    mem[3443] = 8'h00;
    mem[3444] = 8'h00;
    mem[3445] = 8'he0;
    mem[3446] = 8'h00;
    mem[3447] = 8'h07;
    mem[3448] = 8'hf8;
    mem[3449] = 8'h07;
    mem[3450] = 8'h00;
    mem[3451] = 8'h00;
    mem[3452] = 8'h00;
    mem[3453] = 8'h00;
    mem[3454] = 8'h00;
    mem[3455] = 8'h00;
    mem[3456] = 8'h00;
    mem[3457] = 8'h00;
    mem[3458] = 8'h00;
    mem[3459] = 8'h00;
    mem[3460] = 8'hff;
    mem[3461] = 8'h00;
    mem[3462] = 8'hff;
    mem[3463] = 8'h00;
    mem[3464] = 8'h0f;
    mem[3465] = 8'h70;
    mem[3466] = 8'h00;
    mem[3467] = 8'h00;
    mem[3468] = 8'h00;
    mem[3469] = 8'hfe;
    mem[3470] = 8'hff;
    mem[3471] = 8'hff;
    mem[3472] = 8'hff;
    mem[3473] = 8'hff;
    mem[3474] = 8'h0f;
    mem[3475] = 8'h00;
    mem[3476] = 8'h00;
    mem[3477] = 8'he0;
    mem[3478] = 8'h00;
    mem[3479] = 8'h07;
    mem[3480] = 8'hf8;
    mem[3481] = 8'h07;
    mem[3482] = 8'h00;
    mem[3483] = 8'h00;
    mem[3484] = 8'h00;
    mem[3485] = 8'h00;
    mem[3486] = 8'h00;
    mem[3487] = 8'h00;
    mem[3488] = 8'h00;
    mem[3489] = 8'h00;
    mem[3490] = 8'h00;
    mem[3491] = 8'h00;
    mem[3492] = 8'hff;
    mem[3493] = 8'hff;
    mem[3494] = 8'hff;
    mem[3495] = 8'h00;
    mem[3496] = 8'h0f;
    mem[3497] = 8'h70;
    mem[3498] = 8'h00;
    mem[3499] = 8'h00;
    mem[3500] = 8'h00;
    mem[3501] = 8'hfe;
    mem[3502] = 8'hff;
    mem[3503] = 8'hff;
    mem[3504] = 8'hff;
    mem[3505] = 8'hff;
    mem[3506] = 8'h07;
    mem[3507] = 8'h00;
    mem[3508] = 8'h00;
    mem[3509] = 8'he0;
    mem[3510] = 8'h00;
    mem[3511] = 8'h07;
    mem[3512] = 8'hf8;
    mem[3513] = 8'h07;
    mem[3514] = 8'h00;
    mem[3515] = 8'h00;
    mem[3516] = 8'h00;
    mem[3517] = 8'h00;
    mem[3518] = 8'h00;
    mem[3519] = 8'h00;
    mem[3520] = 8'h00;
    mem[3521] = 8'h00;
    mem[3522] = 8'h00;
    mem[3523] = 8'h00;
    mem[3524] = 8'hff;
    mem[3525] = 8'hff;
    mem[3526] = 8'hff;
    mem[3527] = 8'h00;
    mem[3528] = 8'h0f;
    mem[3529] = 8'h70;
    mem[3530] = 8'h00;
    mem[3531] = 8'h00;
    mem[3532] = 8'h00;
    mem[3533] = 8'hfe;
    mem[3534] = 8'hff;
    mem[3535] = 8'hff;
    mem[3536] = 8'hff;
    mem[3537] = 8'hff;
    mem[3538] = 8'h01;
    mem[3539] = 8'h00;
    mem[3540] = 8'h00;
    mem[3541] = 8'he0;
    mem[3542] = 8'h00;
    mem[3543] = 8'h07;
    mem[3544] = 8'hf8;
    mem[3545] = 8'h07;
    mem[3546] = 8'h00;
    mem[3547] = 8'h00;
    mem[3548] = 8'h00;
    mem[3549] = 8'h00;
    mem[3550] = 8'h00;
    mem[3551] = 8'h00;
    mem[3552] = 8'h00;
    mem[3553] = 8'h00;
    mem[3554] = 8'h00;
    mem[3555] = 8'h00;
    mem[3556] = 8'hff;
    mem[3557] = 8'hff;
    mem[3558] = 8'hff;
    mem[3559] = 8'h00;
    mem[3560] = 8'h0f;
    mem[3561] = 8'h70;
    mem[3562] = 8'h00;
    mem[3563] = 8'h00;
    mem[3564] = 8'h00;
    mem[3565] = 8'hfe;
    mem[3566] = 8'hff;
    mem[3567] = 8'hff;
    mem[3568] = 8'hff;
    mem[3569] = 8'hff;
    mem[3570] = 8'h00;
    mem[3571] = 8'h00;
    mem[3572] = 8'h00;
    mem[3573] = 8'he0;
    mem[3574] = 8'h00;
    mem[3575] = 8'h07;
    mem[3576] = 8'hf8;
    mem[3577] = 8'h07;
    mem[3578] = 8'h00;
    mem[3579] = 8'h00;
    mem[3580] = 8'h00;
    mem[3581] = 8'h00;
    mem[3582] = 8'h00;
    mem[3583] = 8'h00;
    mem[3584] = 8'h00;
    mem[3585] = 8'h00;
    mem[3586] = 8'h00;
    mem[3587] = 8'h00;
    mem[3588] = 8'hff;
    mem[3589] = 8'hff;
    mem[3590] = 8'hff;
    mem[3591] = 8'h00;
    mem[3592] = 8'h0f;
    mem[3593] = 8'h70;
    mem[3594] = 8'h00;
    mem[3595] = 8'h00;
    mem[3596] = 8'h00;
    mem[3597] = 8'hfe;
    mem[3598] = 8'hff;
    mem[3599] = 8'hff;
    mem[3600] = 8'hff;
    mem[3601] = 8'hff;
    mem[3602] = 8'h00;
    mem[3603] = 8'h00;
    mem[3604] = 8'h00;
    mem[3605] = 8'he0;
    mem[3606] = 8'h00;
    mem[3607] = 8'h07;
    mem[3608] = 8'hf8;
    mem[3609] = 8'h07;
    mem[3610] = 8'h00;
    mem[3611] = 8'h00;
    mem[3612] = 8'h00;
    mem[3613] = 8'h00;
    mem[3614] = 8'h00;
    mem[3615] = 8'h00;
    mem[3616] = 8'h00;
    mem[3617] = 8'h00;
    mem[3618] = 8'h00;
    mem[3619] = 8'h00;
    mem[3620] = 8'hff;
    mem[3621] = 8'hff;
    mem[3622] = 8'hff;
    mem[3623] = 8'h00;
    mem[3624] = 8'h0f;
    mem[3625] = 8'h70;
    mem[3626] = 8'h00;
    mem[3627] = 8'h00;
    mem[3628] = 8'h00;
    mem[3629] = 8'hfe;
    mem[3630] = 8'hff;
    mem[3631] = 8'hff;
    mem[3632] = 8'hff;
    mem[3633] = 8'hff;
    mem[3634] = 8'h03;
    mem[3635] = 8'h00;
    mem[3636] = 8'h00;
    mem[3637] = 8'he0;
    mem[3638] = 8'h00;
    mem[3639] = 8'h07;
    mem[3640] = 8'hf8;
    mem[3641] = 8'h07;
    mem[3642] = 8'h00;
    mem[3643] = 8'h00;
    mem[3644] = 8'h00;
    mem[3645] = 8'h00;
    mem[3646] = 8'h00;
    mem[3647] = 8'h00;
    mem[3648] = 8'h00;
    mem[3649] = 8'h00;
    mem[3650] = 8'h00;
    mem[3651] = 8'h00;
    mem[3652] = 8'hff;
    mem[3653] = 8'hff;
    mem[3654] = 8'hff;
    mem[3655] = 8'h00;
    mem[3656] = 8'hff;
    mem[3657] = 8'h7f;
    mem[3658] = 8'h00;
    mem[3659] = 8'h00;
    mem[3660] = 8'h00;
    mem[3661] = 8'hfe;
    mem[3662] = 8'hff;
    mem[3663] = 8'hff;
    mem[3664] = 8'hff;
    mem[3665] = 8'hff;
    mem[3666] = 8'h07;
    mem[3667] = 8'h00;
    mem[3668] = 8'h00;
    mem[3669] = 8'he0;
    mem[3670] = 8'h00;
    mem[3671] = 8'h07;
    mem[3672] = 8'hf8;
    mem[3673] = 8'h07;
    mem[3674] = 8'h00;
    mem[3675] = 8'h00;
    mem[3676] = 8'h00;
    mem[3677] = 8'h00;
    mem[3678] = 8'h00;
    mem[3679] = 8'h00;
    mem[3680] = 8'h00;
    mem[3681] = 8'h00;
    mem[3682] = 8'h00;
    mem[3683] = 8'h00;
    mem[3684] = 8'hff;
    mem[3685] = 8'hff;
    mem[3686] = 8'hff;
    mem[3687] = 8'h00;
    mem[3688] = 8'hff;
    mem[3689] = 8'h7f;
    mem[3690] = 8'h00;
    mem[3691] = 8'h00;
    mem[3692] = 8'h00;
    mem[3693] = 8'hfe;
    mem[3694] = 8'hff;
    mem[3695] = 8'hff;
    mem[3696] = 8'hff;
    mem[3697] = 8'hff;
    mem[3698] = 8'h07;
    mem[3699] = 8'h00;
    mem[3700] = 8'h00;
    mem[3701] = 8'he0;
    mem[3702] = 8'h00;
    mem[3703] = 8'h07;
    mem[3704] = 8'hf8;
    mem[3705] = 8'h07;
    mem[3706] = 8'h00;
    mem[3707] = 8'h00;
    mem[3708] = 8'h00;
    mem[3709] = 8'h00;
    mem[3710] = 8'h00;
    mem[3711] = 8'h00;
    mem[3712] = 8'h00;
    mem[3713] = 8'h00;
    mem[3714] = 8'h00;
    mem[3715] = 8'h00;
    mem[3716] = 8'hff;
    mem[3717] = 8'hff;
    mem[3718] = 8'hff;
    mem[3719] = 8'h00;
    mem[3720] = 8'hff;
    mem[3721] = 8'h7f;
    mem[3722] = 8'h00;
    mem[3723] = 8'h00;
    mem[3724] = 8'h00;
    mem[3725] = 8'hfe;
    mem[3726] = 8'hff;
    mem[3727] = 8'hff;
    mem[3728] = 8'hff;
    mem[3729] = 8'hff;
    mem[3730] = 8'h0f;
    mem[3731] = 8'h00;
    mem[3732] = 8'h00;
    mem[3733] = 8'he0;
    mem[3734] = 8'hff;
    mem[3735] = 8'h07;
    mem[3736] = 8'hf8;
    mem[3737] = 8'h07;
    mem[3738] = 8'h00;
    mem[3739] = 8'h00;
    mem[3740] = 8'h00;
    mem[3741] = 8'h00;
    mem[3742] = 8'h00;
    mem[3743] = 8'h00;
    mem[3744] = 8'h00;
    mem[3745] = 8'h00;
    mem[3746] = 8'h00;
    mem[3747] = 8'h00;
    mem[3748] = 8'h00;
    mem[3749] = 8'h00;
    mem[3750] = 8'h00;
    mem[3751] = 8'h00;
    mem[3752] = 8'h0f;
    mem[3753] = 8'h70;
    mem[3754] = 8'h00;
    mem[3755] = 8'h00;
    mem[3756] = 8'h00;
    mem[3757] = 8'hfe;
    mem[3758] = 8'h1f;
    mem[3759] = 8'h00;
    mem[3760] = 8'he0;
    mem[3761] = 8'hff;
    mem[3762] = 8'h0f;
    mem[3763] = 8'h00;
    mem[3764] = 8'h00;
    mem[3765] = 8'he0;
    mem[3766] = 8'hff;
    mem[3767] = 8'h07;
    mem[3768] = 8'h00;
    mem[3769] = 8'h00;
    mem[3770] = 8'hf8;
    mem[3771] = 8'h07;
    mem[3772] = 8'h00;
    mem[3773] = 8'h00;
    mem[3774] = 8'h00;
    mem[3775] = 8'h00;
    mem[3776] = 8'h00;
    mem[3777] = 8'h00;
    mem[3778] = 8'h00;
    mem[3779] = 8'h00;
    mem[3780] = 8'h00;
    mem[3781] = 8'h00;
    mem[3782] = 8'h00;
    mem[3783] = 8'h00;
    mem[3784] = 8'h0f;
    mem[3785] = 8'h70;
    mem[3786] = 8'h00;
    mem[3787] = 8'h00;
    mem[3788] = 8'h00;
    mem[3789] = 8'hfe;
    mem[3790] = 8'h1f;
    mem[3791] = 8'h00;
    mem[3792] = 8'h80;
    mem[3793] = 8'hff;
    mem[3794] = 8'h1f;
    mem[3795] = 8'h00;
    mem[3796] = 8'h00;
    mem[3797] = 8'he0;
    mem[3798] = 8'hff;
    mem[3799] = 8'h07;
    mem[3800] = 8'h00;
    mem[3801] = 8'h00;
    mem[3802] = 8'hf8;
    mem[3803] = 8'h07;
    mem[3804] = 8'h00;
    mem[3805] = 8'h00;
    mem[3806] = 8'h00;
    mem[3807] = 8'h00;
    mem[3808] = 8'h00;
    mem[3809] = 8'h00;
    mem[3810] = 8'h00;
    mem[3811] = 8'h00;
    mem[3812] = 8'h00;
    mem[3813] = 8'h00;
    mem[3814] = 8'h00;
    mem[3815] = 8'h00;
    mem[3816] = 8'h0f;
    mem[3817] = 8'h70;
    mem[3818] = 8'h00;
    mem[3819] = 8'h00;
    mem[3820] = 8'h00;
    mem[3821] = 8'hfe;
    mem[3822] = 8'h1f;
    mem[3823] = 8'h00;
    mem[3824] = 8'h00;
    mem[3825] = 8'hff;
    mem[3826] = 8'h1f;
    mem[3827] = 8'h00;
    mem[3828] = 8'h00;
    mem[3829] = 8'he0;
    mem[3830] = 8'h00;
    mem[3831] = 8'h07;
    mem[3832] = 8'h00;
    mem[3833] = 8'h00;
    mem[3834] = 8'hf8;
    mem[3835] = 8'h07;
    mem[3836] = 8'h00;
    mem[3837] = 8'h00;
    mem[3838] = 8'h00;
    mem[3839] = 8'h00;
    mem[3840] = 8'h00;
    mem[3841] = 8'h00;
    mem[3842] = 8'h00;
    mem[3843] = 8'h00;
    mem[3844] = 8'h00;
    mem[3845] = 8'h00;
    mem[3846] = 8'h00;
    mem[3847] = 8'h00;
    mem[3848] = 8'h0f;
    mem[3849] = 8'h70;
    mem[3850] = 8'h00;
    mem[3851] = 8'h00;
    mem[3852] = 8'h00;
    mem[3853] = 8'hfe;
    mem[3854] = 8'h1f;
    mem[3855] = 8'h00;
    mem[3856] = 8'h00;
    mem[3857] = 8'hfe;
    mem[3858] = 8'h1f;
    mem[3859] = 8'h00;
    mem[3860] = 8'h00;
    mem[3861] = 8'he0;
    mem[3862] = 8'h00;
    mem[3863] = 8'h07;
    mem[3864] = 8'h00;
    mem[3865] = 8'h00;
    mem[3866] = 8'hf8;
    mem[3867] = 8'h07;
    mem[3868] = 8'h00;
    mem[3869] = 8'h00;
    mem[3870] = 8'h00;
    mem[3871] = 8'h00;
    mem[3872] = 8'h00;
    mem[3873] = 8'h00;
    mem[3874] = 8'h00;
    mem[3875] = 8'h00;
    mem[3876] = 8'h00;
    mem[3877] = 8'h00;
    mem[3878] = 8'h00;
    mem[3879] = 8'h00;
    mem[3880] = 8'h0f;
    mem[3881] = 8'h70;
    mem[3882] = 8'h00;
    mem[3883] = 8'h00;
    mem[3884] = 8'h00;
    mem[3885] = 8'hfe;
    mem[3886] = 8'h1f;
    mem[3887] = 8'h00;
    mem[3888] = 8'h00;
    mem[3889] = 8'hfe;
    mem[3890] = 8'h1f;
    mem[3891] = 8'h00;
    mem[3892] = 8'h00;
    mem[3893] = 8'he0;
    mem[3894] = 8'h00;
    mem[3895] = 8'h07;
    mem[3896] = 8'h00;
    mem[3897] = 8'h00;
    mem[3898] = 8'hf8;
    mem[3899] = 8'h07;
    mem[3900] = 8'h00;
    mem[3901] = 8'h00;
    mem[3902] = 8'h00;
    mem[3903] = 8'h00;
    mem[3904] = 8'h00;
    mem[3905] = 8'h00;
    mem[3906] = 8'h00;
    mem[3907] = 8'h00;
    mem[3908] = 8'h00;
    mem[3909] = 8'h00;
    mem[3910] = 8'h00;
    mem[3911] = 8'h00;
    mem[3912] = 8'h0f;
    mem[3913] = 8'h70;
    mem[3914] = 8'h00;
    mem[3915] = 8'h00;
    mem[3916] = 8'h00;
    mem[3917] = 8'hfe;
    mem[3918] = 8'h1f;
    mem[3919] = 8'h00;
    mem[3920] = 8'h00;
    mem[3921] = 8'hfe;
    mem[3922] = 8'h3f;
    mem[3923] = 8'h00;
    mem[3924] = 8'h00;
    mem[3925] = 8'he0;
    mem[3926] = 8'h00;
    mem[3927] = 8'h07;
    mem[3928] = 8'h00;
    mem[3929] = 8'h00;
    mem[3930] = 8'hf8;
    mem[3931] = 8'h07;
    mem[3932] = 8'h00;
    mem[3933] = 8'h00;
    mem[3934] = 8'h00;
    mem[3935] = 8'h00;
    mem[3936] = 8'h00;
    mem[3937] = 8'h00;
    mem[3938] = 8'h00;
    mem[3939] = 8'h00;
    mem[3940] = 8'h00;
    mem[3941] = 8'h00;
    mem[3942] = 8'h00;
    mem[3943] = 8'h00;
    mem[3944] = 8'h0f;
    mem[3945] = 8'h70;
    mem[3946] = 8'h00;
    mem[3947] = 8'h00;
    mem[3948] = 8'h00;
    mem[3949] = 8'hfe;
    mem[3950] = 8'h1f;
    mem[3951] = 8'h00;
    mem[3952] = 8'h00;
    mem[3953] = 8'hfe;
    mem[3954] = 8'h3f;
    mem[3955] = 8'h00;
    mem[3956] = 8'h00;
    mem[3957] = 8'he0;
    mem[3958] = 8'h00;
    mem[3959] = 8'h07;
    mem[3960] = 8'h00;
    mem[3961] = 8'h00;
    mem[3962] = 8'hf8;
    mem[3963] = 8'h07;
    mem[3964] = 8'h00;
    mem[3965] = 8'h00;
    mem[3966] = 8'h00;
    mem[3967] = 8'h00;
    mem[3968] = 8'h00;
    mem[3969] = 8'h00;
    mem[3970] = 8'h00;
    mem[3971] = 8'h00;
    mem[3972] = 8'hff;
    mem[3973] = 8'h00;
    mem[3974] = 8'h00;
    mem[3975] = 8'h00;
    mem[3976] = 8'h0f;
    mem[3977] = 8'h70;
    mem[3978] = 8'h00;
    mem[3979] = 8'h00;
    mem[3980] = 8'h00;
    mem[3981] = 8'hfe;
    mem[3982] = 8'h1f;
    mem[3983] = 8'h00;
    mem[3984] = 8'h00;
    mem[3985] = 8'hfc;
    mem[3986] = 8'h3f;
    mem[3987] = 8'h00;
    mem[3988] = 8'h00;
    mem[3989] = 8'he0;
    mem[3990] = 8'h00;
    mem[3991] = 8'h07;
    mem[3992] = 8'hf8;
    mem[3993] = 8'h07;
    mem[3994] = 8'hf8;
    mem[3995] = 8'h07;
    mem[3996] = 8'h00;
    mem[3997] = 8'h00;
    mem[3998] = 8'h00;
    mem[3999] = 8'h00;
    mem[4000] = 8'h00;
    mem[4001] = 8'h00;
    mem[4002] = 8'h00;
    mem[4003] = 8'h00;
    mem[4004] = 8'hff;
    mem[4005] = 8'h00;
    mem[4006] = 8'hff;
    mem[4007] = 8'h01;
    mem[4008] = 8'h0f;
    mem[4009] = 8'h70;
    mem[4010] = 8'h00;
    mem[4011] = 8'h00;
    mem[4012] = 8'h00;
    mem[4013] = 8'hfe;
    mem[4014] = 8'h1f;
    mem[4015] = 8'h00;
    mem[4016] = 8'h00;
    mem[4017] = 8'hfc;
    mem[4018] = 8'h3f;
    mem[4019] = 8'h00;
    mem[4020] = 8'h00;
    mem[4021] = 8'he0;
    mem[4022] = 8'h00;
    mem[4023] = 8'h07;
    mem[4024] = 8'hf8;
    mem[4025] = 8'h07;
    mem[4026] = 8'hf8;
    mem[4027] = 8'h07;
    mem[4028] = 8'h00;
    mem[4029] = 8'h00;
    mem[4030] = 8'h00;
    mem[4031] = 8'h00;
    mem[4032] = 8'h00;
    mem[4033] = 8'h00;
    mem[4034] = 8'h00;
    mem[4035] = 8'h00;
    mem[4036] = 8'hff;
    mem[4037] = 8'h80;
    mem[4038] = 8'hff;
    mem[4039] = 8'h03;
    mem[4040] = 8'h0f;
    mem[4041] = 8'h70;
    mem[4042] = 8'h00;
    mem[4043] = 8'h00;
    mem[4044] = 8'h00;
    mem[4045] = 8'hfe;
    mem[4046] = 8'h1f;
    mem[4047] = 8'h00;
    mem[4048] = 8'h00;
    mem[4049] = 8'hfc;
    mem[4050] = 8'h3f;
    mem[4051] = 8'h00;
    mem[4052] = 8'h00;
    mem[4053] = 8'he0;
    mem[4054] = 8'h00;
    mem[4055] = 8'h07;
    mem[4056] = 8'hf8;
    mem[4057] = 8'h07;
    mem[4058] = 8'hf8;
    mem[4059] = 8'h07;
    mem[4060] = 8'h00;
    mem[4061] = 8'h00;
    mem[4062] = 8'h00;
    mem[4063] = 8'h00;
    mem[4064] = 8'h00;
    mem[4065] = 8'h00;
    mem[4066] = 8'h00;
    mem[4067] = 8'h00;
    mem[4068] = 8'hff;
    mem[4069] = 8'hc0;
    mem[4070] = 8'hff;
    mem[4071] = 8'h07;
    mem[4072] = 8'h0f;
    mem[4073] = 8'h70;
    mem[4074] = 8'h00;
    mem[4075] = 8'h00;
    mem[4076] = 8'h00;
    mem[4077] = 8'hfe;
    mem[4078] = 8'h1f;
    mem[4079] = 8'h00;
    mem[4080] = 8'h00;
    mem[4081] = 8'hfc;
    mem[4082] = 8'h3f;
    mem[4083] = 8'h00;
    mem[4084] = 8'h00;
    mem[4085] = 8'he0;
    mem[4086] = 8'h00;
    mem[4087] = 8'h07;
    mem[4088] = 8'hf8;
    mem[4089] = 8'h07;
    mem[4090] = 8'hf8;
    mem[4091] = 8'h07;
    mem[4092] = 8'h00;
    mem[4093] = 8'h00;
    mem[4094] = 8'h00;
    mem[4095] = 8'h00;
    mem[4096] = 8'h00;
    mem[4097] = 8'h00;
    mem[4098] = 8'h00;
    mem[4099] = 8'h00;
    mem[4100] = 8'hff;
    mem[4101] = 8'he0;
    mem[4102] = 8'hff;
    mem[4103] = 8'h0f;
    mem[4104] = 8'h0f;
    mem[4105] = 8'h70;
    mem[4106] = 8'h00;
    mem[4107] = 8'h00;
    mem[4108] = 8'h00;
    mem[4109] = 8'hfe;
    mem[4110] = 8'h1f;
    mem[4111] = 8'h00;
    mem[4112] = 8'h00;
    mem[4113] = 8'hfc;
    mem[4114] = 8'h3f;
    mem[4115] = 8'h00;
    mem[4116] = 8'h00;
    mem[4117] = 8'he0;
    mem[4118] = 8'h00;
    mem[4119] = 8'h07;
    mem[4120] = 8'hf8;
    mem[4121] = 8'h07;
    mem[4122] = 8'hf8;
    mem[4123] = 8'h07;
    mem[4124] = 8'h00;
    mem[4125] = 8'h00;
    mem[4126] = 8'h00;
    mem[4127] = 8'h00;
    mem[4128] = 8'h00;
    mem[4129] = 8'h00;
    mem[4130] = 8'h00;
    mem[4131] = 8'h00;
    mem[4132] = 8'hff;
    mem[4133] = 8'he0;
    mem[4134] = 8'hc7;
    mem[4135] = 8'h0f;
    mem[4136] = 8'h0f;
    mem[4137] = 8'h70;
    mem[4138] = 8'h00;
    mem[4139] = 8'h00;
    mem[4140] = 8'h00;
    mem[4141] = 8'hfe;
    mem[4142] = 8'h1f;
    mem[4143] = 8'h00;
    mem[4144] = 8'h00;
    mem[4145] = 8'hfc;
    mem[4146] = 8'h3f;
    mem[4147] = 8'h00;
    mem[4148] = 8'h00;
    mem[4149] = 8'he0;
    mem[4150] = 8'h00;
    mem[4151] = 8'h07;
    mem[4152] = 8'hf8;
    mem[4153] = 8'h07;
    mem[4154] = 8'hf8;
    mem[4155] = 8'h07;
    mem[4156] = 8'h00;
    mem[4157] = 8'h00;
    mem[4158] = 8'h00;
    mem[4159] = 8'h00;
    mem[4160] = 8'h00;
    mem[4161] = 8'h00;
    mem[4162] = 8'h00;
    mem[4163] = 8'h00;
    mem[4164] = 8'hff;
    mem[4165] = 8'hf0;
    mem[4166] = 8'h83;
    mem[4167] = 8'h1f;
    mem[4168] = 8'h0f;
    mem[4169] = 8'h70;
    mem[4170] = 8'h00;
    mem[4171] = 8'h00;
    mem[4172] = 8'h00;
    mem[4173] = 8'hfe;
    mem[4174] = 8'h1f;
    mem[4175] = 8'h00;
    mem[4176] = 8'h00;
    mem[4177] = 8'hfc;
    mem[4178] = 8'h3f;
    mem[4179] = 8'h00;
    mem[4180] = 8'h00;
    mem[4181] = 8'he0;
    mem[4182] = 8'h00;
    mem[4183] = 8'h07;
    mem[4184] = 8'hf8;
    mem[4185] = 8'h07;
    mem[4186] = 8'hf8;
    mem[4187] = 8'h07;
    mem[4188] = 8'h00;
    mem[4189] = 8'h00;
    mem[4190] = 8'h00;
    mem[4191] = 8'h00;
    mem[4192] = 8'h00;
    mem[4193] = 8'h00;
    mem[4194] = 8'h00;
    mem[4195] = 8'h00;
    mem[4196] = 8'hff;
    mem[4197] = 8'hf0;
    mem[4198] = 8'h01;
    mem[4199] = 8'h1f;
    mem[4200] = 8'h0f;
    mem[4201] = 8'h70;
    mem[4202] = 8'h00;
    mem[4203] = 8'h00;
    mem[4204] = 8'h00;
    mem[4205] = 8'hfe;
    mem[4206] = 8'h1f;
    mem[4207] = 8'h00;
    mem[4208] = 8'h00;
    mem[4209] = 8'hfc;
    mem[4210] = 8'h3f;
    mem[4211] = 8'h00;
    mem[4212] = 8'h00;
    mem[4213] = 8'he0;
    mem[4214] = 8'h00;
    mem[4215] = 8'h07;
    mem[4216] = 8'hf8;
    mem[4217] = 8'h07;
    mem[4218] = 8'hf8;
    mem[4219] = 8'h07;
    mem[4220] = 8'h00;
    mem[4221] = 8'h00;
    mem[4222] = 8'h00;
    mem[4223] = 8'h00;
    mem[4224] = 8'h00;
    mem[4225] = 8'h00;
    mem[4226] = 8'h00;
    mem[4227] = 8'h00;
    mem[4228] = 8'hff;
    mem[4229] = 8'hf0;
    mem[4230] = 8'h01;
    mem[4231] = 8'h1f;
    mem[4232] = 8'h0f;
    mem[4233] = 8'h70;
    mem[4234] = 8'h00;
    mem[4235] = 8'h00;
    mem[4236] = 8'h00;
    mem[4237] = 8'hfe;
    mem[4238] = 8'h1f;
    mem[4239] = 8'h00;
    mem[4240] = 8'h00;
    mem[4241] = 8'hfc;
    mem[4242] = 8'h3f;
    mem[4243] = 8'h00;
    mem[4244] = 8'h00;
    mem[4245] = 8'he0;
    mem[4246] = 8'h00;
    mem[4247] = 8'h07;
    mem[4248] = 8'hf8;
    mem[4249] = 8'h07;
    mem[4250] = 8'hf8;
    mem[4251] = 8'h07;
    mem[4252] = 8'h00;
    mem[4253] = 8'h00;
    mem[4254] = 8'h00;
    mem[4255] = 8'h00;
    mem[4256] = 8'h00;
    mem[4257] = 8'h00;
    mem[4258] = 8'h00;
    mem[4259] = 8'h00;
    mem[4260] = 8'hff;
    mem[4261] = 8'hf0;
    mem[4262] = 8'h00;
    mem[4263] = 8'h1e;
    mem[4264] = 8'h0f;
    mem[4265] = 8'h70;
    mem[4266] = 8'h00;
    mem[4267] = 8'h00;
    mem[4268] = 8'h00;
    mem[4269] = 8'hfe;
    mem[4270] = 8'h1f;
    mem[4271] = 8'h00;
    mem[4272] = 8'h00;
    mem[4273] = 8'hfc;
    mem[4274] = 8'h3f;
    mem[4275] = 8'h00;
    mem[4276] = 8'h00;
    mem[4277] = 8'he0;
    mem[4278] = 8'h00;
    mem[4279] = 8'h07;
    mem[4280] = 8'hf8;
    mem[4281] = 8'h07;
    mem[4282] = 8'hf8;
    mem[4283] = 8'h07;
    mem[4284] = 8'h00;
    mem[4285] = 8'h00;
    mem[4286] = 8'h00;
    mem[4287] = 8'h00;
    mem[4288] = 8'h00;
    mem[4289] = 8'h00;
    mem[4290] = 8'h00;
    mem[4291] = 8'h00;
    mem[4292] = 8'hff;
    mem[4293] = 8'hf0;
    mem[4294] = 8'h01;
    mem[4295] = 8'h1f;
    mem[4296] = 8'h0f;
    mem[4297] = 8'h70;
    mem[4298] = 8'h00;
    mem[4299] = 8'h00;
    mem[4300] = 8'h00;
    mem[4301] = 8'hfe;
    mem[4302] = 8'h1f;
    mem[4303] = 8'h00;
    mem[4304] = 8'h00;
    mem[4305] = 8'hfc;
    mem[4306] = 8'h3f;
    mem[4307] = 8'h00;
    mem[4308] = 8'h00;
    mem[4309] = 8'he0;
    mem[4310] = 8'h00;
    mem[4311] = 8'h07;
    mem[4312] = 8'hf8;
    mem[4313] = 8'h07;
    mem[4314] = 8'hf8;
    mem[4315] = 8'h07;
    mem[4316] = 8'h00;
    mem[4317] = 8'h00;
    mem[4318] = 8'h00;
    mem[4319] = 8'h00;
    mem[4320] = 8'h00;
    mem[4321] = 8'h00;
    mem[4322] = 8'h00;
    mem[4323] = 8'h00;
    mem[4324] = 8'hfe;
    mem[4325] = 8'hf0;
    mem[4326] = 8'h01;
    mem[4327] = 8'h1f;
    mem[4328] = 8'h0f;
    mem[4329] = 8'h70;
    mem[4330] = 8'h00;
    mem[4331] = 8'h00;
    mem[4332] = 8'h00;
    mem[4333] = 8'hfe;
    mem[4334] = 8'h1f;
    mem[4335] = 8'h00;
    mem[4336] = 8'h00;
    mem[4337] = 8'hfc;
    mem[4338] = 8'h3f;
    mem[4339] = 8'h00;
    mem[4340] = 8'h00;
    mem[4341] = 8'he0;
    mem[4342] = 8'h00;
    mem[4343] = 8'h07;
    mem[4344] = 8'hf8;
    mem[4345] = 8'h07;
    mem[4346] = 8'hf8;
    mem[4347] = 8'h07;
    mem[4348] = 8'h00;
    mem[4349] = 8'h00;
    mem[4350] = 8'h00;
    mem[4351] = 8'h00;
    mem[4352] = 8'h00;
    mem[4353] = 8'h00;
    mem[4354] = 8'h00;
    mem[4355] = 8'h00;
    mem[4356] = 8'hfe;
    mem[4357] = 8'hf0;
    mem[4358] = 8'h83;
    mem[4359] = 8'h1f;
    mem[4360] = 8'h0f;
    mem[4361] = 8'h70;
    mem[4362] = 8'h00;
    mem[4363] = 8'h00;
    mem[4364] = 8'h00;
    mem[4365] = 8'hfe;
    mem[4366] = 8'h1f;
    mem[4367] = 8'h00;
    mem[4368] = 8'h00;
    mem[4369] = 8'hfc;
    mem[4370] = 8'h3f;
    mem[4371] = 8'h00;
    mem[4372] = 8'h00;
    mem[4373] = 8'he0;
    mem[4374] = 8'h00;
    mem[4375] = 8'h07;
    mem[4376] = 8'hf8;
    mem[4377] = 8'h07;
    mem[4378] = 8'hf8;
    mem[4379] = 8'h07;
    mem[4380] = 8'h00;
    mem[4381] = 8'h00;
    mem[4382] = 8'h00;
    mem[4383] = 8'h00;
    mem[4384] = 8'h00;
    mem[4385] = 8'h00;
    mem[4386] = 8'h00;
    mem[4387] = 8'h00;
    mem[4388] = 8'hfe;
    mem[4389] = 8'he0;
    mem[4390] = 8'hff;
    mem[4391] = 8'h0f;
    mem[4392] = 8'h0f;
    mem[4393] = 8'h70;
    mem[4394] = 8'h00;
    mem[4395] = 8'h00;
    mem[4396] = 8'h00;
    mem[4397] = 8'hfe;
    mem[4398] = 8'h1f;
    mem[4399] = 8'h00;
    mem[4400] = 8'h00;
    mem[4401] = 8'hfc;
    mem[4402] = 8'h7f;
    mem[4403] = 8'h00;
    mem[4404] = 8'h00;
    mem[4405] = 8'he0;
    mem[4406] = 8'h00;
    mem[4407] = 8'h07;
    mem[4408] = 8'hf8;
    mem[4409] = 8'h07;
    mem[4410] = 8'hf8;
    mem[4411] = 8'h07;
    mem[4412] = 8'h00;
    mem[4413] = 8'h00;
    mem[4414] = 8'h00;
    mem[4415] = 8'h00;
    mem[4416] = 8'h00;
    mem[4417] = 8'h00;
    mem[4418] = 8'h00;
    mem[4419] = 8'h00;
    mem[4420] = 8'hfe;
    mem[4421] = 8'hc0;
    mem[4422] = 8'hff;
    mem[4423] = 8'h07;
    mem[4424] = 8'h0f;
    mem[4425] = 8'h70;
    mem[4426] = 8'h00;
    mem[4427] = 8'h00;
    mem[4428] = 8'h00;
    mem[4429] = 8'hfe;
    mem[4430] = 8'h1f;
    mem[4431] = 8'h00;
    mem[4432] = 8'h00;
    mem[4433] = 8'hf8;
    mem[4434] = 8'h7f;
    mem[4435] = 8'h00;
    mem[4436] = 8'h00;
    mem[4437] = 8'he0;
    mem[4438] = 8'h00;
    mem[4439] = 8'h07;
    mem[4440] = 8'hf8;
    mem[4441] = 8'h07;
    mem[4442] = 8'hf8;
    mem[4443] = 8'h07;
    mem[4444] = 8'h00;
    mem[4445] = 8'h00;
    mem[4446] = 8'h00;
    mem[4447] = 8'h00;
    mem[4448] = 8'h00;
    mem[4449] = 8'h00;
    mem[4450] = 8'h00;
    mem[4451] = 8'h00;
    mem[4452] = 8'hfe;
    mem[4453] = 8'h80;
    mem[4454] = 8'hff;
    mem[4455] = 8'h07;
    mem[4456] = 8'h0f;
    mem[4457] = 8'h70;
    mem[4458] = 8'h00;
    mem[4459] = 8'h00;
    mem[4460] = 8'h00;
    mem[4461] = 8'hfe;
    mem[4462] = 8'h1f;
    mem[4463] = 8'h00;
    mem[4464] = 8'h00;
    mem[4465] = 8'hf8;
    mem[4466] = 8'h7f;
    mem[4467] = 8'h00;
    mem[4468] = 8'h00;
    mem[4469] = 8'he0;
    mem[4470] = 8'h7e;
    mem[4471] = 8'h07;
    mem[4472] = 8'hf8;
    mem[4473] = 8'h07;
    mem[4474] = 8'hf8;
    mem[4475] = 8'h07;
    mem[4476] = 8'h00;
    mem[4477] = 8'h00;
    mem[4478] = 8'h00;
    mem[4479] = 8'h00;
    mem[4480] = 8'h00;
    mem[4481] = 8'h00;
    mem[4482] = 8'h00;
    mem[4483] = 8'h00;
    mem[4484] = 8'hfe;
    mem[4485] = 8'h00;
    mem[4486] = 8'hff;
    mem[4487] = 8'h01;
    mem[4488] = 8'h0f;
    mem[4489] = 8'h70;
    mem[4490] = 8'h00;
    mem[4491] = 8'h00;
    mem[4492] = 8'h00;
    mem[4493] = 8'h00;
    mem[4494] = 8'h00;
    mem[4495] = 8'h00;
    mem[4496] = 8'h00;
    mem[4497] = 8'h00;
    mem[4498] = 8'h00;
    mem[4499] = 8'h00;
    mem[4500] = 8'h00;
    mem[4501] = 8'he0;
    mem[4502] = 8'hff;
    mem[4503] = 8'h07;
    mem[4504] = 8'hf8;
    mem[4505] = 8'h07;
    mem[4506] = 8'hf8;
    mem[4507] = 8'h07;
    mem[4508] = 8'h00;
    mem[4509] = 8'h00;
    mem[4510] = 8'h00;
    mem[4511] = 8'h00;
    mem[4512] = 8'h00;
    mem[4513] = 8'h00;
    mem[4514] = 8'h00;
    mem[4515] = 8'h00;
    mem[4516] = 8'hfe;
    mem[4517] = 8'h00;
    mem[4518] = 8'hfe;
    mem[4519] = 8'h01;
    mem[4520] = 8'h0f;
    mem[4521] = 8'h70;
    mem[4522] = 8'h00;
    mem[4523] = 8'h00;
    mem[4524] = 8'h00;
    mem[4525] = 8'hfe;
    mem[4526] = 8'hff;
    mem[4527] = 8'hff;
    mem[4528] = 8'hff;
    mem[4529] = 8'hff;
    mem[4530] = 8'h7f;
    mem[4531] = 8'h00;
    mem[4532] = 8'h00;
    mem[4533] = 8'he0;
    mem[4534] = 8'hff;
    mem[4535] = 8'h07;
    mem[4536] = 8'hf8;
    mem[4537] = 8'h07;
    mem[4538] = 8'hf8;
    mem[4539] = 8'h07;
    mem[4540] = 8'h00;
    mem[4541] = 8'h00;
    mem[4542] = 8'h00;
    mem[4543] = 8'h00;
    mem[4544] = 8'h00;
    mem[4545] = 8'h00;
    mem[4546] = 8'h00;
    mem[4547] = 8'h00;
    mem[4548] = 8'hfe;
    mem[4549] = 8'h00;
    mem[4550] = 8'hfe;
    mem[4551] = 8'h01;
    mem[4552] = 8'h0f;
    mem[4553] = 8'h70;
    mem[4554] = 8'h00;
    mem[4555] = 8'h00;
    mem[4556] = 8'h00;
    mem[4557] = 8'h00;
    mem[4558] = 8'h00;
    mem[4559] = 8'h00;
    mem[4560] = 8'h00;
    mem[4561] = 8'h00;
    mem[4562] = 8'h00;
    mem[4563] = 8'h00;
    mem[4564] = 8'h00;
    mem[4565] = 8'he0;
    mem[4566] = 8'hc3;
    mem[4567] = 8'h07;
    mem[4568] = 8'hf8;
    mem[4569] = 8'h03;
    mem[4570] = 8'hf8;
    mem[4571] = 8'h07;
    mem[4572] = 8'h00;
    mem[4573] = 8'h00;
    mem[4574] = 8'h00;
    mem[4575] = 8'h00;
    mem[4576] = 8'h00;
    mem[4577] = 8'h00;
    mem[4578] = 8'h00;
    mem[4579] = 8'h00;
    mem[4580] = 8'hfe;
    mem[4581] = 8'h00;
    mem[4582] = 8'hfe;
    mem[4583] = 8'h01;
    mem[4584] = 8'h1e;
    mem[4585] = 8'h70;
    mem[4586] = 8'h00;
    mem[4587] = 8'h00;
    mem[4588] = 8'h00;
    mem[4589] = 8'h00;
    mem[4590] = 8'h00;
    mem[4591] = 8'h00;
    mem[4592] = 8'h00;
    mem[4593] = 8'h00;
    mem[4594] = 8'h00;
    mem[4595] = 8'h00;
    mem[4596] = 8'h00;
    mem[4597] = 8'he0;
    mem[4598] = 8'h00;
    mem[4599] = 8'h07;
    mem[4600] = 8'hf8;
    mem[4601] = 8'h03;
    mem[4602] = 8'hf8;
    mem[4603] = 8'h07;
    mem[4604] = 8'h00;
    mem[4605] = 8'h00;
    mem[4606] = 8'h00;
    mem[4607] = 8'h00;
    mem[4608] = 8'h00;
    mem[4609] = 8'h00;
    mem[4610] = 8'h00;
    mem[4611] = 8'h00;
    mem[4612] = 8'hfe;
    mem[4613] = 8'h00;
    mem[4614] = 8'hfe;
    mem[4615] = 8'h01;
    mem[4616] = 8'h3e;
    mem[4617] = 8'h70;
    mem[4618] = 8'h00;
    mem[4619] = 8'h00;
    mem[4620] = 8'h00;
    mem[4621] = 8'h00;
    mem[4622] = 8'h00;
    mem[4623] = 8'h00;
    mem[4624] = 8'h00;
    mem[4625] = 8'h00;
    mem[4626] = 8'h00;
    mem[4627] = 8'h00;
    mem[4628] = 8'h00;
    mem[4629] = 8'h70;
    mem[4630] = 8'h7e;
    mem[4631] = 8'h0e;
    mem[4632] = 8'hf8;
    mem[4633] = 8'h03;
    mem[4634] = 8'hf8;
    mem[4635] = 8'h07;
    mem[4636] = 8'h00;
    mem[4637] = 8'h00;
    mem[4638] = 8'h00;
    mem[4639] = 8'h00;
    mem[4640] = 8'h00;
    mem[4641] = 8'h00;
    mem[4642] = 8'h00;
    mem[4643] = 8'h00;
    mem[4644] = 8'hfe;
    mem[4645] = 8'h00;
    mem[4646] = 8'hfe;
    mem[4647] = 8'h01;
    mem[4648] = 8'hfe;
    mem[4649] = 8'h70;
    mem[4650] = 8'h00;
    mem[4651] = 8'h00;
    mem[4652] = 8'h00;
    mem[4653] = 8'h00;
    mem[4654] = 8'h3c;
    mem[4655] = 8'h8f;
    mem[4656] = 8'hf7;
    mem[4657] = 8'h3d;
    mem[4658] = 8'h00;
    mem[4659] = 8'h00;
    mem[4660] = 8'h00;
    mem[4661] = 8'h70;
    mem[4662] = 8'h7e;
    mem[4663] = 8'h0e;
    mem[4664] = 8'hf8;
    mem[4665] = 8'h03;
    mem[4666] = 8'hf8;
    mem[4667] = 8'h07;
    mem[4668] = 8'h00;
    mem[4669] = 8'h00;
    mem[4670] = 8'h00;
    mem[4671] = 8'h00;
    mem[4672] = 8'h00;
    mem[4673] = 8'h00;
    mem[4674] = 8'h00;
    mem[4675] = 8'h00;
    mem[4676] = 8'hfe;
    mem[4677] = 8'h01;
    mem[4678] = 8'hfe;
    mem[4679] = 8'h01;
    mem[4680] = 8'hfe;
    mem[4681] = 8'h71;
    mem[4682] = 8'h00;
    mem[4683] = 8'h00;
    mem[4684] = 8'h00;
    mem[4685] = 8'h00;
    mem[4686] = 8'h64;
    mem[4687] = 8'hd1;
    mem[4688] = 8'h4c;
    mem[4689] = 8'h04;
    mem[4690] = 8'h00;
    mem[4691] = 8'h00;
    mem[4692] = 8'h00;
    mem[4693] = 8'h7c;
    mem[4694] = 8'hff;
    mem[4695] = 8'h0e;
    mem[4696] = 8'hf8;
    mem[4697] = 8'h03;
    mem[4698] = 8'hf8;
    mem[4699] = 8'h07;
    mem[4700] = 8'h00;
    mem[4701] = 8'h00;
    mem[4702] = 8'h00;
    mem[4703] = 8'h00;
    mem[4704] = 8'h00;
    mem[4705] = 8'h00;
    mem[4706] = 8'h00;
    mem[4707] = 8'h00;
    mem[4708] = 8'hfe;
    mem[4709] = 8'h01;
    mem[4710] = 8'hfe;
    mem[4711] = 8'h01;
    mem[4712] = 8'hfe;
    mem[4713] = 8'h77;
    mem[4714] = 8'h00;
    mem[4715] = 8'h00;
    mem[4716] = 8'h00;
    mem[4717] = 8'h00;
    mem[4718] = 8'ha4;
    mem[4719] = 8'hd1;
    mem[4720] = 8'h48;
    mem[4721] = 8'h0c;
    mem[4722] = 8'h00;
    mem[4723] = 8'h00;
    mem[4724] = 8'h00;
    mem[4725] = 8'h7e;
    mem[4726] = 8'he7;
    mem[4727] = 8'h0e;
    mem[4728] = 8'hf8;
    mem[4729] = 8'h03;
    mem[4730] = 8'hf8;
    mem[4731] = 8'h07;
    mem[4732] = 8'h00;
    mem[4733] = 8'h00;
    mem[4734] = 8'h00;
    mem[4735] = 8'h00;
    mem[4736] = 8'h00;
    mem[4737] = 8'h00;
    mem[4738] = 8'h00;
    mem[4739] = 8'h00;
    mem[4740] = 8'hfe;
    mem[4741] = 8'h01;
    mem[4742] = 8'hfe;
    mem[4743] = 8'h01;
    mem[4744] = 8'hfe;
    mem[4745] = 8'h7f;
    mem[4746] = 8'h00;
    mem[4747] = 8'h00;
    mem[4748] = 8'h00;
    mem[4749] = 8'h00;
    mem[4750] = 8'h9c;
    mem[4751] = 8'hd1;
    mem[4752] = 8'h48;
    mem[4753] = 8'h38;
    mem[4754] = 8'h00;
    mem[4755] = 8'h00;
    mem[4756] = 8'h80;
    mem[4757] = 8'h7f;
    mem[4758] = 8'hff;
    mem[4759] = 8'h0e;
    mem[4760] = 8'hf8;
    mem[4761] = 8'h03;
    mem[4762] = 8'hf8;
    mem[4763] = 8'h03;
    mem[4764] = 8'h00;
    mem[4765] = 8'h00;
    mem[4766] = 8'h00;
    mem[4767] = 8'h00;
    mem[4768] = 8'h00;
    mem[4769] = 8'h00;
    mem[4770] = 8'h00;
    mem[4771] = 8'h00;
    mem[4772] = 8'hfe;
    mem[4773] = 8'h01;
    mem[4774] = 8'hfe;
    mem[4775] = 8'h01;
    mem[4776] = 8'hfc;
    mem[4777] = 8'h7f;
    mem[4778] = 8'h00;
    mem[4779] = 8'h00;
    mem[4780] = 8'h00;
    mem[4781] = 8'h00;
    mem[4782] = 8'h24;
    mem[4783] = 8'hd9;
    mem[4784] = 8'h4c;
    mem[4785] = 8'h30;
    mem[4786] = 8'h00;
    mem[4787] = 8'h00;
    mem[4788] = 8'hc0;
    mem[4789] = 8'h77;
    mem[4790] = 8'hff;
    mem[4791] = 8'h0e;
    mem[4792] = 8'hf8;
    mem[4793] = 8'h03;
    mem[4794] = 8'hf8;
    mem[4795] = 8'h03;
    mem[4796] = 8'h00;
    mem[4797] = 8'h00;
    mem[4798] = 8'h00;
    mem[4799] = 8'h00;
    mem[4800] = 8'h00;
    mem[4801] = 8'h00;
    mem[4802] = 8'h00;
    mem[4803] = 8'h00;
    mem[4804] = 8'hfe;
    mem[4805] = 8'h01;
    mem[4806] = 8'hfe;
    mem[4807] = 8'h01;
    mem[4808] = 8'hf8;
    mem[4809] = 8'hff;
    mem[4810] = 8'h00;
    mem[4811] = 8'h00;
    mem[4812] = 8'h00;
    mem[4813] = 8'h00;
    mem[4814] = 8'h64;
    mem[4815] = 8'h8f;
    mem[4816] = 8'h47;
    mem[4817] = 8'h1c;
    mem[4818] = 8'h00;
    mem[4819] = 8'h00;
    mem[4820] = 8'hf0;
    mem[4821] = 8'h73;
    mem[4822] = 8'h7e;
    mem[4823] = 8'h0e;
    mem[4824] = 8'hfc;
    mem[4825] = 8'h03;
    mem[4826] = 8'hf8;
    mem[4827] = 8'h03;
    mem[4828] = 8'h00;
    mem[4829] = 8'h00;
    mem[4830] = 8'h00;
    mem[4831] = 8'h00;
    mem[4832] = 8'h00;
    mem[4833] = 8'h00;
    mem[4834] = 8'h00;
    mem[4835] = 8'h00;
    mem[4836] = 8'hfe;
    mem[4837] = 8'h01;
    mem[4838] = 8'hfc;
    mem[4839] = 8'h01;
    mem[4840] = 8'hf0;
    mem[4841] = 8'hff;
    mem[4842] = 8'h03;
    mem[4843] = 8'h00;
    mem[4844] = 8'h00;
    mem[4845] = 8'h00;
    mem[4846] = 8'h00;
    mem[4847] = 8'h00;
    mem[4848] = 8'h00;
    mem[4849] = 8'h00;
    mem[4850] = 8'h00;
    mem[4851] = 8'h00;
    mem[4852] = 8'hf8;
    mem[4853] = 8'he0;
    mem[4854] = 8'h18;
    mem[4855] = 8'h07;
    mem[4856] = 8'hfc;
    mem[4857] = 8'h03;
    mem[4858] = 8'hf8;
    mem[4859] = 8'h03;
    mem[4860] = 8'h00;
    mem[4861] = 8'h00;
    mem[4862] = 8'h00;
    mem[4863] = 8'h00;
    mem[4864] = 8'h00;
    mem[4865] = 8'h00;
    mem[4866] = 8'h00;
    mem[4867] = 8'h00;
    mem[4868] = 8'hfe;
    mem[4869] = 8'h01;
    mem[4870] = 8'hfc;
    mem[4871] = 8'h01;
    mem[4872] = 8'he0;
    mem[4873] = 8'hff;
    mem[4874] = 8'h07;
    mem[4875] = 8'h00;
    mem[4876] = 8'h00;
    mem[4877] = 8'h00;
    mem[4878] = 8'h00;
    mem[4879] = 8'h00;
    mem[4880] = 8'h00;
    mem[4881] = 8'h00;
    mem[4882] = 8'h00;
    mem[4883] = 8'h00;
    mem[4884] = 8'h7e;
    mem[4885] = 8'he0;
    mem[4886] = 8'hc3;
    mem[4887] = 8'h07;
    mem[4888] = 8'hfc;
    mem[4889] = 8'h03;
    mem[4890] = 8'hf8;
    mem[4891] = 8'h03;
    mem[4892] = 8'h00;
    mem[4893] = 8'h00;
    mem[4894] = 8'h00;
    mem[4895] = 8'h00;
    mem[4896] = 8'h00;
    mem[4897] = 8'h00;
    mem[4898] = 8'h00;
    mem[4899] = 8'h00;
    mem[4900] = 8'hfe;
    mem[4901] = 8'h01;
    mem[4902] = 8'hfc;
    mem[4903] = 8'h01;
    mem[4904] = 8'hc0;
    mem[4905] = 8'hff;
    mem[4906] = 8'h1f;
    mem[4907] = 8'h00;
    mem[4908] = 8'h00;
    mem[4909] = 8'h00;
    mem[4910] = 8'h00;
    mem[4911] = 8'h00;
    mem[4912] = 8'h00;
    mem[4913] = 8'h00;
    mem[4914] = 8'h00;
    mem[4915] = 8'h00;
    mem[4916] = 8'h1f;
    mem[4917] = 8'hc0;
    mem[4918] = 8'hff;
    mem[4919] = 8'h03;
    mem[4920] = 8'hfc;
    mem[4921] = 8'h03;
    mem[4922] = 8'hf8;
    mem[4923] = 8'h03;
    mem[4924] = 8'h00;
    mem[4925] = 8'h00;
    mem[4926] = 8'h00;
    mem[4927] = 8'h00;
    mem[4928] = 8'h00;
    mem[4929] = 8'h00;
    mem[4930] = 8'h00;
    mem[4931] = 8'h00;
    mem[4932] = 8'hfe;
    mem[4933] = 8'h01;
    mem[4934] = 8'hfc;
    mem[4935] = 8'h01;
    mem[4936] = 8'h80;
    mem[4937] = 8'hff;
    mem[4938] = 8'h7f;
    mem[4939] = 8'h00;
    mem[4940] = 8'h00;
    mem[4941] = 8'h00;
    mem[4942] = 8'h00;
    mem[4943] = 8'h70;
    mem[4944] = 8'h00;
    mem[4945] = 8'h00;
    mem[4946] = 8'h00;
    mem[4947] = 8'hc0;
    mem[4948] = 8'h0f;
    mem[4949] = 8'h80;
    mem[4950] = 8'hff;
    mem[4951] = 8'h01;
    mem[4952] = 8'hfc;
    mem[4953] = 8'h03;
    mem[4954] = 8'hf8;
    mem[4955] = 8'h03;
    mem[4956] = 8'h00;
    mem[4957] = 8'h00;
    mem[4958] = 8'h00;
    mem[4959] = 8'h00;
    mem[4960] = 8'h00;
    mem[4961] = 8'h00;
    mem[4962] = 8'h00;
    mem[4963] = 8'h00;
    mem[4964] = 8'hfe;
    mem[4965] = 8'h01;
    mem[4966] = 8'hfc;
    mem[4967] = 8'h03;
    mem[4968] = 8'h00;
    mem[4969] = 8'hfe;
    mem[4970] = 8'hff;
    mem[4971] = 8'h01;
    mem[4972] = 8'h00;
    mem[4973] = 8'h00;
    mem[4974] = 8'h00;
    mem[4975] = 8'h70;
    mem[4976] = 8'h00;
    mem[4977] = 8'h00;
    mem[4978] = 8'h00;
    mem[4979] = 8'he0;
    mem[4980] = 8'h03;
    mem[4981] = 8'h80;
    mem[4982] = 8'h7f;
    mem[4983] = 8'h00;
    mem[4984] = 8'hfc;
    mem[4985] = 8'h01;
    mem[4986] = 8'hfc;
    mem[4987] = 8'h03;
    mem[4988] = 8'h00;
    mem[4989] = 8'h00;
    mem[4990] = 8'h00;
    mem[4991] = 8'h00;
    mem[4992] = 8'h00;
    mem[4993] = 8'h00;
    mem[4994] = 8'h00;
    mem[4995] = 8'h00;
    mem[4996] = 8'hfe;
    mem[4997] = 8'h01;
    mem[4998] = 8'hfc;
    mem[4999] = 8'h03;
    mem[5000] = 8'h00;
    mem[5001] = 8'hfc;
    mem[5002] = 8'hff;
    mem[5003] = 8'h03;
    mem[5004] = 8'h00;
    mem[5005] = 8'h00;
    mem[5006] = 8'h00;
    mem[5007] = 8'h70;
    mem[5008] = 8'h00;
    mem[5009] = 8'h00;
    mem[5010] = 8'h80;
    mem[5011] = 8'hff;
    mem[5012] = 8'h01;
    mem[5013] = 8'he0;
    mem[5014] = 8'h07;
    mem[5015] = 8'h00;
    mem[5016] = 8'hfe;
    mem[5017] = 8'h01;
    mem[5018] = 8'hfc;
    mem[5019] = 8'h03;
    mem[5020] = 8'h00;
    mem[5021] = 8'h00;
    mem[5022] = 8'h00;
    mem[5023] = 8'h00;
    mem[5024] = 8'h00;
    mem[5025] = 8'h00;
    mem[5026] = 8'h00;
    mem[5027] = 8'h00;
    mem[5028] = 8'hfe;
    mem[5029] = 8'h01;
    mem[5030] = 8'hfc;
    mem[5031] = 8'h0f;
    mem[5032] = 8'h00;
    mem[5033] = 8'hf0;
    mem[5034] = 8'hff;
    mem[5035] = 8'h0f;
    mem[5036] = 8'h00;
    mem[5037] = 8'h00;
    mem[5038] = 8'h00;
    mem[5039] = 8'h70;
    mem[5040] = 8'h00;
    mem[5041] = 8'h00;
    mem[5042] = 8'he0;
    mem[5043] = 8'h7f;
    mem[5044] = 8'h00;
    mem[5045] = 8'hf0;
    mem[5046] = 8'h01;
    mem[5047] = 8'h00;
    mem[5048] = 8'hff;
    mem[5049] = 8'h01;
    mem[5050] = 8'hfc;
    mem[5051] = 8'h03;
    mem[5052] = 8'h00;
    mem[5053] = 8'h00;
    mem[5054] = 8'h00;
    mem[5055] = 8'h00;
    mem[5056] = 8'h00;
    mem[5057] = 8'h00;
    mem[5058] = 8'h00;
    mem[5059] = 8'h00;
    mem[5060] = 8'hfc;
    mem[5061] = 8'h01;
    mem[5062] = 8'hfc;
    mem[5063] = 8'h1f;
    mem[5064] = 8'h00;
    mem[5065] = 8'he0;
    mem[5066] = 8'hff;
    mem[5067] = 8'h9f;
    mem[5068] = 8'h0f;
    mem[5069] = 8'h00;
    mem[5070] = 8'h00;
    mem[5071] = 8'h70;
    mem[5072] = 8'h00;
    mem[5073] = 8'h00;
    mem[5074] = 8'hf0;
    mem[5075] = 8'hff;
    mem[5076] = 8'h01;
    mem[5077] = 8'hfc;
    mem[5078] = 8'h00;
    mem[5079] = 8'hc0;
    mem[5080] = 8'hff;
    mem[5081] = 8'h01;
    mem[5082] = 8'hfc;
    mem[5083] = 8'h03;
    mem[5084] = 8'h00;
    mem[5085] = 8'h00;
    mem[5086] = 8'h00;
    mem[5087] = 8'h00;
    mem[5088] = 8'h00;
    mem[5089] = 8'h00;
    mem[5090] = 8'h00;
    mem[5091] = 8'h00;
    mem[5092] = 8'hfc;
    mem[5093] = 8'h01;
    mem[5094] = 8'hf8;
    mem[5095] = 8'h3f;
    mem[5096] = 8'h00;
    mem[5097] = 8'h80;
    mem[5098] = 8'hff;
    mem[5099] = 8'hff;
    mem[5100] = 8'h7f;
    mem[5101] = 8'h00;
    mem[5102] = 8'h00;
    mem[5103] = 8'hfe;
    mem[5104] = 8'h03;
    mem[5105] = 8'h00;
    mem[5106] = 8'hf0;
    mem[5107] = 8'he0;
    mem[5108] = 8'h01;
    mem[5109] = 8'h3f;
    mem[5110] = 8'h00;
    mem[5111] = 8'he0;
    mem[5112] = 8'hff;
    mem[5113] = 8'h00;
    mem[5114] = 8'hfc;
    mem[5115] = 8'h03;
    mem[5116] = 8'h00;
    mem[5117] = 8'h00;
    mem[5118] = 8'h00;
    mem[5119] = 8'h00;
    mem[5120] = 8'h00;
    mem[5121] = 8'h00;
    mem[5122] = 8'h00;
    mem[5123] = 8'h00;
    mem[5124] = 8'hfc;
    mem[5125] = 8'h01;
    mem[5126] = 8'hf0;
    mem[5127] = 8'hff;
    mem[5128] = 8'h00;
    mem[5129] = 8'h00;
    mem[5130] = 8'hff;
    mem[5131] = 8'hff;
    mem[5132] = 8'hff;
    mem[5133] = 8'h00;
    mem[5134] = 8'h00;
    mem[5135] = 8'hfe;
    mem[5136] = 8'h03;
    mem[5137] = 8'h00;
    mem[5138] = 8'h78;
    mem[5139] = 8'hce;
    mem[5140] = 8'h83;
    mem[5141] = 8'h1f;
    mem[5142] = 8'h00;
    mem[5143] = 8'hf8;
    mem[5144] = 8'hff;
    mem[5145] = 8'h00;
    mem[5146] = 8'hfc;
    mem[5147] = 8'h03;
    mem[5148] = 8'h00;
    mem[5149] = 8'h00;
    mem[5150] = 8'h00;
    mem[5151] = 8'h00;
    mem[5152] = 8'h00;
    mem[5153] = 8'h00;
    mem[5154] = 8'h00;
    mem[5155] = 8'h00;
    mem[5156] = 8'hfc;
    mem[5157] = 8'h01;
    mem[5158] = 8'he0;
    mem[5159] = 8'hff;
    mem[5160] = 8'h01;
    mem[5161] = 8'h00;
    mem[5162] = 8'hfc;
    mem[5163] = 8'hff;
    mem[5164] = 8'hff;
    mem[5165] = 8'h01;
    mem[5166] = 8'h00;
    mem[5167] = 8'hfe;
    mem[5168] = 8'h03;
    mem[5169] = 8'h00;
    mem[5170] = 8'h3c;
    mem[5171] = 8'h9f;
    mem[5172] = 8'he3;
    mem[5173] = 8'h07;
    mem[5174] = 8'h00;
    mem[5175] = 8'hfc;
    mem[5176] = 8'h7f;
    mem[5177] = 8'h00;
    mem[5178] = 8'hfc;
    mem[5179] = 8'h03;
    mem[5180] = 8'h00;
    mem[5181] = 8'h00;
    mem[5182] = 8'h00;
    mem[5183] = 8'h00;
    mem[5184] = 8'h00;
    mem[5185] = 8'h00;
    mem[5186] = 8'h00;
    mem[5187] = 8'h00;
    mem[5188] = 8'hfc;
    mem[5189] = 8'h03;
    mem[5190] = 8'hc0;
    mem[5191] = 8'hff;
    mem[5192] = 8'h07;
    mem[5193] = 8'h00;
    mem[5194] = 8'hf0;
    mem[5195] = 8'hff;
    mem[5196] = 8'hff;
    mem[5197] = 8'h01;
    mem[5198] = 8'h00;
    mem[5199] = 8'h8e;
    mem[5200] = 8'h03;
    mem[5201] = 8'h00;
    mem[5202] = 8'h9f;
    mem[5203] = 8'h3f;
    mem[5204] = 8'hf7;
    mem[5205] = 8'h01;
    mem[5206] = 8'h00;
    mem[5207] = 8'hff;
    mem[5208] = 8'h1f;
    mem[5209] = 8'h00;
    mem[5210] = 8'hfc;
    mem[5211] = 8'h01;
    mem[5212] = 8'h00;
    mem[5213] = 8'h00;
    mem[5214] = 8'h00;
    mem[5215] = 8'h00;
    mem[5216] = 8'h00;
    mem[5217] = 8'h00;
    mem[5218] = 8'h00;
    mem[5219] = 8'h00;
    mem[5220] = 8'hfc;
    mem[5221] = 8'h03;
    mem[5222] = 8'h80;
    mem[5223] = 8'hff;
    mem[5224] = 8'h1f;
    mem[5225] = 8'h00;
    mem[5226] = 8'he0;
    mem[5227] = 8'h7f;
    mem[5228] = 8'hf0;
    mem[5229] = 8'h03;
    mem[5230] = 8'h80;
    mem[5231] = 8'hff;
    mem[5232] = 8'h0f;
    mem[5233] = 8'hc0;
    mem[5234] = 8'hdf;
    mem[5235] = 8'h3b;
    mem[5236] = 8'hff;
    mem[5237] = 8'h00;
    mem[5238] = 8'hc0;
    mem[5239] = 8'hff;
    mem[5240] = 8'h0f;
    mem[5241] = 8'h00;
    mem[5242] = 8'hfc;
    mem[5243] = 8'h01;
    mem[5244] = 8'h00;
    mem[5245] = 8'h00;
    mem[5246] = 8'h00;
    mem[5247] = 8'h00;
    mem[5248] = 8'h00;
    mem[5249] = 8'h00;
    mem[5250] = 8'h00;
    mem[5251] = 8'h00;
    mem[5252] = 8'hfc;
    mem[5253] = 8'h03;
    mem[5254] = 8'h00;
    mem[5255] = 8'hfe;
    mem[5256] = 8'h3f;
    mem[5257] = 8'h00;
    mem[5258] = 8'h80;
    mem[5259] = 8'h3f;
    mem[5260] = 8'he0;
    mem[5261] = 8'h03;
    mem[5262] = 8'h80;
    mem[5263] = 8'hff;
    mem[5264] = 8'h0f;
    mem[5265] = 8'hf0;
    mem[5266] = 8'hdf;
    mem[5267] = 8'h39;
    mem[5268] = 8'h3f;
    mem[5269] = 8'h00;
    mem[5270] = 8'he0;
    mem[5271] = 8'hff;
    mem[5272] = 8'h07;
    mem[5273] = 8'h00;
    mem[5274] = 8'hfe;
    mem[5275] = 8'h01;
    mem[5276] = 8'h00;
    mem[5277] = 8'h00;
    mem[5278] = 8'h00;
    mem[5279] = 8'h00;
    mem[5280] = 8'h00;
    mem[5281] = 8'h00;
    mem[5282] = 8'h00;
    mem[5283] = 8'h00;
    mem[5284] = 8'hfc;
    mem[5285] = 8'h07;
    mem[5286] = 8'h00;
    mem[5287] = 8'hfc;
    mem[5288] = 8'hff;
    mem[5289] = 8'h00;
    mem[5290] = 8'h00;
    mem[5291] = 8'h3f;
    mem[5292] = 8'he0;
    mem[5293] = 8'h03;
    mem[5294] = 8'h80;
    mem[5295] = 8'hff;
    mem[5296] = 8'h0f;
    mem[5297] = 8'hf8;
    mem[5298] = 8'h9d;
    mem[5299] = 8'h3f;
    mem[5300] = 8'h1f;
    mem[5301] = 8'h00;
    mem[5302] = 8'hf8;
    mem[5303] = 8'hff;
    mem[5304] = 8'h01;
    mem[5305] = 8'h00;
    mem[5306] = 8'hfe;
    mem[5307] = 8'h01;
    mem[5308] = 8'h00;
    mem[5309] = 8'h00;
    mem[5310] = 8'h00;
    mem[5311] = 8'h00;
    mem[5312] = 8'h00;
    mem[5313] = 8'h00;
    mem[5314] = 8'h00;
    mem[5315] = 8'h00;
    mem[5316] = 8'hf8;
    mem[5317] = 8'h0f;
    mem[5318] = 8'h00;
    mem[5319] = 8'hf0;
    mem[5320] = 8'hff;
    mem[5321] = 8'h01;
    mem[5322] = 8'h00;
    mem[5323] = 8'h3e;
    mem[5324] = 8'hc0;
    mem[5325] = 8'h03;
    mem[5326] = 8'h80;
    mem[5327] = 8'h73;
    mem[5328] = 8'h0e;
    mem[5329] = 8'h7e;
    mem[5330] = 8'h9c;
    mem[5331] = 8'hbf;
    mem[5332] = 8'h07;
    mem[5333] = 8'h00;
    mem[5334] = 8'hfc;
    mem[5335] = 8'hff;
    mem[5336] = 8'h00;
    mem[5337] = 8'h00;
    mem[5338] = 8'hff;
    mem[5339] = 8'h01;
    mem[5340] = 8'h00;
    mem[5341] = 8'h00;
    mem[5342] = 8'h00;
    mem[5343] = 8'h00;
    mem[5344] = 8'h00;
    mem[5345] = 8'h00;
    mem[5346] = 8'h00;
    mem[5347] = 8'h00;
    mem[5348] = 8'hf8;
    mem[5349] = 8'h1f;
    mem[5350] = 8'h00;
    mem[5351] = 8'he0;
    mem[5352] = 8'hff;
    mem[5353] = 8'h07;
    mem[5354] = 8'h00;
    mem[5355] = 8'h3e;
    mem[5356] = 8'hc0;
    mem[5357] = 8'h03;
    mem[5358] = 8'h80;
    mem[5359] = 8'h73;
    mem[5360] = 8'h8e;
    mem[5361] = 8'h1f;
    mem[5362] = 8'h38;
    mem[5363] = 8'h9f;
    mem[5364] = 8'h03;
    mem[5365] = 8'h00;
    mem[5366] = 8'hff;
    mem[5367] = 8'h3f;
    mem[5368] = 8'h00;
    mem[5369] = 8'hc0;
    mem[5370] = 8'hff;
    mem[5371] = 8'h01;
    mem[5372] = 8'h00;
    mem[5373] = 8'h00;
    mem[5374] = 8'h00;
    mem[5375] = 8'h00;
    mem[5376] = 8'h00;
    mem[5377] = 8'h00;
    mem[5378] = 8'h00;
    mem[5379] = 8'h00;
    mem[5380] = 8'hf8;
    mem[5381] = 8'h7f;
    mem[5382] = 8'h00;
    mem[5383] = 8'hc0;
    mem[5384] = 8'hff;
    mem[5385] = 8'h1f;
    mem[5386] = 8'h00;
    mem[5387] = 8'h3e;
    mem[5388] = 8'he0;
    mem[5389] = 8'h03;
    mem[5390] = 8'h80;
    mem[5391] = 8'h73;
    mem[5392] = 8'hee;
    mem[5393] = 8'h07;
    mem[5394] = 8'h78;
    mem[5395] = 8'hc0;
    mem[5396] = 8'h03;
    mem[5397] = 8'hc0;
    mem[5398] = 8'hff;
    mem[5399] = 8'h1f;
    mem[5400] = 8'h00;
    mem[5401] = 8'he0;
    mem[5402] = 8'hff;
    mem[5403] = 8'h00;
    mem[5404] = 8'h00;
    mem[5405] = 8'h00;
    mem[5406] = 8'h00;
    mem[5407] = 8'h00;
    mem[5408] = 8'h00;
    mem[5409] = 8'h00;
    mem[5410] = 8'h00;
    mem[5411] = 8'h00;
    mem[5412] = 8'hf0;
    mem[5413] = 8'hff;
    mem[5414] = 8'h00;
    mem[5415] = 8'h00;
    mem[5416] = 8'hff;
    mem[5417] = 8'h3f;
    mem[5418] = 8'h00;
    mem[5419] = 8'h7e;
    mem[5420] = 8'he0;
    mem[5421] = 8'h03;
    mem[5422] = 8'h80;
    mem[5423] = 8'h73;
    mem[5424] = 8'hfe;
    mem[5425] = 8'h03;
    mem[5426] = 8'hf0;
    mem[5427] = 8'hf1;
    mem[5428] = 8'h01;
    mem[5429] = 8'he0;
    mem[5430] = 8'hff;
    mem[5431] = 8'h07;
    mem[5432] = 8'h00;
    mem[5433] = 8'hf8;
    mem[5434] = 8'hff;
    mem[5435] = 8'h00;
    mem[5436] = 8'h00;
    mem[5437] = 8'h00;
    mem[5438] = 8'h00;
    mem[5439] = 8'h00;
    mem[5440] = 8'h00;
    mem[5441] = 8'h00;
    mem[5442] = 8'h00;
    mem[5443] = 8'h00;
    mem[5444] = 8'he0;
    mem[5445] = 8'hff;
    mem[5446] = 8'h03;
    mem[5447] = 8'h00;
    mem[5448] = 8'hfc;
    mem[5449] = 8'hff;
    mem[5450] = 8'h00;
    mem[5451] = 8'hfc;
    mem[5452] = 8'hf8;
    mem[5453] = 8'h01;
    mem[5454] = 8'h80;
    mem[5455] = 8'h73;
    mem[5456] = 8'hfe;
    mem[5457] = 8'h00;
    mem[5458] = 8'he0;
    mem[5459] = 8'hff;
    mem[5460] = 8'h00;
    mem[5461] = 8'hf8;
    mem[5462] = 8'hff;
    mem[5463] = 8'h03;
    mem[5464] = 8'h00;
    mem[5465] = 8'hfc;
    mem[5466] = 8'h7f;
    mem[5467] = 8'h00;
    mem[5468] = 8'h00;
    mem[5469] = 8'h00;
    mem[5470] = 8'h00;
    mem[5471] = 8'h00;
    mem[5472] = 8'h00;
    mem[5473] = 8'h00;
    mem[5474] = 8'h00;
    mem[5475] = 8'h00;
    mem[5476] = 8'hc0;
    mem[5477] = 8'hff;
    mem[5478] = 8'h07;
    mem[5479] = 8'h00;
    mem[5480] = 8'hf8;
    mem[5481] = 8'hff;
    mem[5482] = 8'h03;
    mem[5483] = 8'hfc;
    mem[5484] = 8'hff;
    mem[5485] = 8'h01;
    mem[5486] = 8'h80;
    mem[5487] = 8'hff;
    mem[5488] = 8'h3f;
    mem[5489] = 8'h00;
    mem[5490] = 8'hf0;
    mem[5491] = 8'h7f;
    mem[5492] = 8'h00;
    mem[5493] = 8'hfe;
    mem[5494] = 8'hff;
    mem[5495] = 8'h00;
    mem[5496] = 8'h00;
    mem[5497] = 8'hff;
    mem[5498] = 8'h1f;
    mem[5499] = 8'h00;
    mem[5500] = 8'h00;
    mem[5501] = 8'h00;
    mem[5502] = 8'h00;
    mem[5503] = 8'h00;
    mem[5504] = 8'h00;
    mem[5505] = 8'h00;
    mem[5506] = 8'h00;
    mem[5507] = 8'h00;
    mem[5508] = 8'h80;
    mem[5509] = 8'hff;
    mem[5510] = 8'h1f;
    mem[5511] = 8'h00;
    mem[5512] = 8'he0;
    mem[5513] = 8'hff;
    mem[5514] = 8'h07;
    mem[5515] = 8'hf8;
    mem[5516] = 8'hff;
    mem[5517] = 8'h00;
    mem[5518] = 8'h80;
    mem[5519] = 8'hff;
    mem[5520] = 8'h0f;
    mem[5521] = 8'h00;
    mem[5522] = 8'hfc;
    mem[5523] = 8'h1f;
    mem[5524] = 8'h00;
    mem[5525] = 8'hff;
    mem[5526] = 8'h7f;
    mem[5527] = 8'h00;
    mem[5528] = 8'h80;
    mem[5529] = 8'hff;
    mem[5530] = 8'h0f;
    mem[5531] = 8'h00;
    mem[5532] = 8'h00;
    mem[5533] = 8'h00;
    mem[5534] = 8'h00;
    mem[5535] = 8'h00;
    mem[5536] = 8'h00;
    mem[5537] = 8'h00;
    mem[5538] = 8'h00;
    mem[5539] = 8'h00;
    mem[5540] = 8'h00;
    mem[5541] = 8'hfe;
    mem[5542] = 8'h3f;
    mem[5543] = 8'h7f;
    mem[5544] = 8'hc0;
    mem[5545] = 8'hff;
    mem[5546] = 8'h1f;
    mem[5547] = 8'hf0;
    mem[5548] = 8'h7f;
    mem[5549] = 8'h00;
    mem[5550] = 8'h80;
    mem[5551] = 8'hff;
    mem[5552] = 8'h0f;
    mem[5553] = 8'h00;
    mem[5554] = 8'h3f;
    mem[5555] = 8'h00;
    mem[5556] = 8'hc0;
    mem[5557] = 8'hff;
    mem[5558] = 8'h1f;
    mem[5559] = 8'h00;
    mem[5560] = 8'he0;
    mem[5561] = 8'hff;
    mem[5562] = 8'h07;
    mem[5563] = 8'h00;
    mem[5564] = 8'h00;
    mem[5565] = 8'h00;
    mem[5566] = 8'h00;
    mem[5567] = 8'h00;
    mem[5568] = 8'h00;
    mem[5569] = 8'h00;
    mem[5570] = 8'h00;
    mem[5571] = 8'h00;
    mem[5572] = 8'h00;
    mem[5573] = 8'hfc;
    mem[5574] = 8'hff;
    mem[5575] = 8'hff;
    mem[5576] = 8'h01;
    mem[5577] = 8'hff;
    mem[5578] = 8'h7f;
    mem[5579] = 8'hc0;
    mem[5580] = 8'h3f;
    mem[5581] = 8'h00;
    mem[5582] = 8'h80;
    mem[5583] = 8'h07;
    mem[5584] = 8'h1f;
    mem[5585] = 8'h80;
    mem[5586] = 8'h1f;
    mem[5587] = 8'h00;
    mem[5588] = 8'hf0;
    mem[5589] = 8'hff;
    mem[5590] = 8'h07;
    mem[5591] = 8'h00;
    mem[5592] = 8'hf0;
    mem[5593] = 8'hff;
    mem[5594] = 8'h01;
    mem[5595] = 8'h00;
    mem[5596] = 8'h00;
    mem[5597] = 8'h00;
    mem[5598] = 8'h00;
    mem[5599] = 8'h00;
    mem[5600] = 8'h00;
    mem[5601] = 8'h00;
    mem[5602] = 8'h00;
    mem[5603] = 8'h00;
    mem[5604] = 8'h00;
    mem[5605] = 8'hf0;
    mem[5606] = 8'hff;
    mem[5607] = 8'hff;
    mem[5608] = 8'h03;
    mem[5609] = 8'hfc;
    mem[5610] = 8'hff;
    mem[5611] = 8'h01;
    mem[5612] = 8'h00;
    mem[5613] = 8'h00;
    mem[5614] = 8'hc0;
    mem[5615] = 8'h73;
    mem[5616] = 8'h1c;
    mem[5617] = 8'he0;
    mem[5618] = 8'h07;
    mem[5619] = 8'h00;
    mem[5620] = 8'hf8;
    mem[5621] = 8'hff;
    mem[5622] = 8'h03;
    mem[5623] = 8'h00;
    mem[5624] = 8'hfc;
    mem[5625] = 8'hff;
    mem[5626] = 8'h00;
    mem[5627] = 8'h00;
    mem[5628] = 8'h00;
    mem[5629] = 8'h00;
    mem[5630] = 8'h00;
    mem[5631] = 8'h00;
    mem[5632] = 8'h00;
    mem[5633] = 8'h00;
    mem[5634] = 8'h00;
    mem[5635] = 8'h00;
    mem[5636] = 8'h00;
    mem[5637] = 8'he0;
    mem[5638] = 8'hff;
    mem[5639] = 8'hff;
    mem[5640] = 8'h07;
    mem[5641] = 8'hf8;
    mem[5642] = 8'hff;
    mem[5643] = 8'h03;
    mem[5644] = 8'h00;
    mem[5645] = 8'h00;
    mem[5646] = 8'hc0;
    mem[5647] = 8'hf9;
    mem[5648] = 8'h3d;
    mem[5649] = 8'hf8;
    mem[5650] = 8'h01;
    mem[5651] = 8'h00;
    mem[5652] = 8'hfe;
    mem[5653] = 8'hff;
    mem[5654] = 8'h00;
    mem[5655] = 8'h00;
    mem[5656] = 8'hff;
    mem[5657] = 8'h7f;
    mem[5658] = 8'h00;
    mem[5659] = 8'h00;
    mem[5660] = 8'h00;
    mem[5661] = 8'h00;
    mem[5662] = 8'h00;
    mem[5663] = 8'h00;
    mem[5664] = 8'h00;
    mem[5665] = 8'h00;
    mem[5666] = 8'h00;
    mem[5667] = 8'h00;
    mem[5668] = 8'h00;
    mem[5669] = 8'h80;
    mem[5670] = 8'hff;
    mem[5671] = 8'hf7;
    mem[5672] = 8'h07;
    mem[5673] = 8'he0;
    mem[5674] = 8'hff;
    mem[5675] = 8'h0f;
    mem[5676] = 8'h00;
    mem[5677] = 8'h00;
    mem[5678] = 8'he0;
    mem[5679] = 8'hfd;
    mem[5680] = 8'h39;
    mem[5681] = 8'h7e;
    mem[5682] = 8'h00;
    mem[5683] = 8'h80;
    mem[5684] = 8'hff;
    mem[5685] = 8'h7f;
    mem[5686] = 8'h00;
    mem[5687] = 8'h80;
    mem[5688] = 8'hff;
    mem[5689] = 8'h1f;
    mem[5690] = 8'h00;
    mem[5691] = 8'h00;
    mem[5692] = 8'h00;
    mem[5693] = 8'h00;
    mem[5694] = 8'h00;
    mem[5695] = 8'h00;
    mem[5696] = 8'h00;
    mem[5697] = 8'h00;
    mem[5698] = 8'h00;
    mem[5699] = 8'h00;
    mem[5700] = 8'h00;
    mem[5701] = 8'h00;
    mem[5702] = 8'hff;
    mem[5703] = 8'hc1;
    mem[5704] = 8'h0f;
    mem[5705] = 8'h80;
    mem[5706] = 8'hff;
    mem[5707] = 8'h3f;
    mem[5708] = 8'h00;
    mem[5709] = 8'h00;
    mem[5710] = 8'he0;
    mem[5711] = 8'hdc;
    mem[5712] = 8'hbb;
    mem[5713] = 8'h3f;
    mem[5714] = 8'h00;
    mem[5715] = 8'he0;
    mem[5716] = 8'hff;
    mem[5717] = 8'h1f;
    mem[5718] = 8'h00;
    mem[5719] = 8'he0;
    mem[5720] = 8'hff;
    mem[5721] = 8'h07;
    mem[5722] = 8'h00;
    mem[5723] = 8'h00;
    mem[5724] = 8'h00;
    mem[5725] = 8'h00;
    mem[5726] = 8'h00;
    mem[5727] = 8'h00;
    mem[5728] = 8'h00;
    mem[5729] = 8'h00;
    mem[5730] = 8'h00;
    mem[5731] = 8'h00;
    mem[5732] = 8'h00;
    mem[5733] = 8'h00;
    mem[5734] = 8'hfc;
    mem[5735] = 8'h80;
    mem[5736] = 8'h0f;
    mem[5737] = 8'h00;
    mem[5738] = 8'hff;
    mem[5739] = 8'hff;
    mem[5740] = 8'h00;
    mem[5741] = 8'h00;
    mem[5742] = 8'he0;
    mem[5743] = 8'h9c;
    mem[5744] = 8'hfb;
    mem[5745] = 8'h0f;
    mem[5746] = 8'h00;
    mem[5747] = 8'hf0;
    mem[5748] = 8'hff;
    mem[5749] = 8'h07;
    mem[5750] = 8'h00;
    mem[5751] = 8'hf8;
    mem[5752] = 8'hff;
    mem[5753] = 8'h03;
    mem[5754] = 8'h00;
    mem[5755] = 8'h00;
    mem[5756] = 8'h00;
    mem[5757] = 8'h00;
    mem[5758] = 8'h00;
    mem[5759] = 8'h00;
    mem[5760] = 8'h00;
    mem[5761] = 8'h00;
    mem[5762] = 8'h00;
    mem[5763] = 8'h00;
    mem[5764] = 8'h00;
    mem[5765] = 8'h00;
    mem[5766] = 8'hf8;
    mem[5767] = 8'h00;
    mem[5768] = 8'h0f;
    mem[5769] = 8'h00;
    mem[5770] = 8'hfc;
    mem[5771] = 8'hff;
    mem[5772] = 8'h01;
    mem[5773] = 8'h00;
    mem[5774] = 8'he0;
    mem[5775] = 8'hfc;
    mem[5776] = 8'hfb;
    mem[5777] = 8'h03;
    mem[5778] = 8'h00;
    mem[5779] = 8'hfc;
    mem[5780] = 8'hff;
    mem[5781] = 8'h01;
    mem[5782] = 8'h00;
    mem[5783] = 8'hfc;
    mem[5784] = 8'hff;
    mem[5785] = 8'h00;
    mem[5786] = 8'h00;
    mem[5787] = 8'h00;
    mem[5788] = 8'h00;
    mem[5789] = 8'h00;
    mem[5790] = 8'h00;
    mem[5791] = 8'h00;
    mem[5792] = 8'h00;
    mem[5793] = 8'h00;
    mem[5794] = 8'h00;
    mem[5795] = 8'h00;
    mem[5796] = 8'h00;
    mem[5797] = 8'h00;
    mem[5798] = 8'hf8;
    mem[5799] = 8'h00;
    mem[5800] = 8'h0f;
    mem[5801] = 8'h00;
    mem[5802] = 8'hf0;
    mem[5803] = 8'hff;
    mem[5804] = 8'h07;
    mem[5805] = 8'h00;
    mem[5806] = 8'hc0;
    mem[5807] = 8'hfd;
    mem[5808] = 8'hf9;
    mem[5809] = 8'h00;
    mem[5810] = 8'h00;
    mem[5811] = 8'hff;
    mem[5812] = 8'hff;
    mem[5813] = 8'h00;
    mem[5814] = 8'h00;
    mem[5815] = 8'hff;
    mem[5816] = 8'h7f;
    mem[5817] = 8'h00;
    mem[5818] = 8'h00;
    mem[5819] = 8'h00;
    mem[5820] = 8'h00;
    mem[5821] = 8'h00;
    mem[5822] = 8'h00;
    mem[5823] = 8'h00;
    mem[5824] = 8'h00;
    mem[5825] = 8'h00;
    mem[5826] = 8'h00;
    mem[5827] = 8'h00;
    mem[5828] = 8'h00;
    mem[5829] = 8'h00;
    mem[5830] = 8'hf8;
    mem[5831] = 8'h00;
    mem[5832] = 8'h0f;
    mem[5833] = 8'h00;
    mem[5834] = 8'he0;
    mem[5835] = 8'hff;
    mem[5836] = 8'h1f;
    mem[5837] = 8'h00;
    mem[5838] = 8'hc0;
    mem[5839] = 8'hf9;
    mem[5840] = 8'h7c;
    mem[5841] = 8'h00;
    mem[5842] = 8'h80;
    mem[5843] = 8'hff;
    mem[5844] = 8'h3f;
    mem[5845] = 8'h00;
    mem[5846] = 8'hc0;
    mem[5847] = 8'hff;
    mem[5848] = 8'h1f;
    mem[5849] = 8'h00;
    mem[5850] = 8'h00;
    mem[5851] = 8'h00;
    mem[5852] = 8'h00;
    mem[5853] = 8'h00;
    mem[5854] = 8'h00;
    mem[5855] = 8'h00;
    mem[5856] = 8'h00;
    mem[5857] = 8'h00;
    mem[5858] = 8'h00;
    mem[5859] = 8'h00;
    mem[5860] = 8'h00;
    mem[5861] = 8'h00;
    mem[5862] = 8'hf8;
    mem[5863] = 8'h80;
    mem[5864] = 8'h0f;
    mem[5865] = 8'h00;
    mem[5866] = 8'h80;
    mem[5867] = 8'hff;
    mem[5868] = 8'h7f;
    mem[5869] = 8'h00;
    mem[5870] = 8'hc0;
    mem[5871] = 8'h03;
    mem[5872] = 8'h1e;
    mem[5873] = 8'h00;
    mem[5874] = 8'h80;
    mem[5875] = 8'hff;
    mem[5876] = 8'h1f;
    mem[5877] = 8'h00;
    mem[5878] = 8'he0;
    mem[5879] = 8'hff;
    mem[5880] = 8'h0f;
    mem[5881] = 8'h00;
    mem[5882] = 8'h00;
    mem[5883] = 8'h00;
    mem[5884] = 8'h00;
    mem[5885] = 8'h00;
    mem[5886] = 8'h00;
    mem[5887] = 8'h00;
    mem[5888] = 8'h00;
    mem[5889] = 8'h00;
    mem[5890] = 8'h00;
    mem[5891] = 8'h00;
    mem[5892] = 8'h00;
    mem[5893] = 8'h00;
    mem[5894] = 8'hf8;
    mem[5895] = 8'hc1;
    mem[5896] = 8'h0f;
    mem[5897] = 8'h00;
    mem[5898] = 8'h00;
    mem[5899] = 8'hfe;
    mem[5900] = 8'hff;
    mem[5901] = 8'h01;
    mem[5902] = 8'h80;
    mem[5903] = 8'h8f;
    mem[5904] = 8'h0f;
    mem[5905] = 8'h00;
    mem[5906] = 8'h80;
    mem[5907] = 8'hff;
    mem[5908] = 8'h07;
    mem[5909] = 8'h00;
    mem[5910] = 8'hf8;
    mem[5911] = 8'hff;
    mem[5912] = 8'h03;
    mem[5913] = 8'h00;
    mem[5914] = 8'h00;
    mem[5915] = 8'h00;
    mem[5916] = 8'h00;
    mem[5917] = 8'h00;
    mem[5918] = 8'h00;
    mem[5919] = 8'h00;
    mem[5920] = 8'h00;
    mem[5921] = 8'h00;
    mem[5922] = 8'h00;
    mem[5923] = 8'h00;
    mem[5924] = 8'h00;
    mem[5925] = 8'h00;
    mem[5926] = 8'hf0;
    mem[5927] = 8'hf7;
    mem[5928] = 8'h07;
    mem[5929] = 8'h00;
    mem[5930] = 8'h00;
    mem[5931] = 8'hf8;
    mem[5932] = 8'hff;
    mem[5933] = 8'h03;
    mem[5934] = 8'h00;
    mem[5935] = 8'hff;
    mem[5936] = 8'h07;
    mem[5937] = 8'h00;
    mem[5938] = 8'h00;
    mem[5939] = 8'hff;
    mem[5940] = 8'h01;
    mem[5941] = 8'h00;
    mem[5942] = 8'hfe;
    mem[5943] = 8'hff;
    mem[5944] = 8'h01;
    mem[5945] = 8'h00;
    mem[5946] = 8'h00;
    mem[5947] = 8'h00;
    mem[5948] = 8'h00;
    mem[5949] = 8'h00;
    mem[5950] = 8'h00;
    mem[5951] = 8'h00;
    mem[5952] = 8'h00;
    mem[5953] = 8'h00;
    mem[5954] = 8'h00;
    mem[5955] = 8'h00;
    mem[5956] = 8'h00;
    mem[5957] = 8'h00;
    mem[5958] = 8'he0;
    mem[5959] = 8'hff;
    mem[5960] = 8'h07;
    mem[5961] = 8'h00;
    mem[5962] = 8'h00;
    mem[5963] = 8'hf0;
    mem[5964] = 8'hff;
    mem[5965] = 8'h0f;
    mem[5966] = 8'h00;
    mem[5967] = 8'hfe;
    mem[5968] = 8'h03;
    mem[5969] = 8'h80;
    mem[5970] = 8'h03;
    mem[5971] = 8'h7e;
    mem[5972] = 8'h00;
    mem[5973] = 8'h00;
    mem[5974] = 8'hff;
    mem[5975] = 8'h7f;
    mem[5976] = 8'h00;
    mem[5977] = 8'h00;
    mem[5978] = 8'h00;
    mem[5979] = 8'h00;
    mem[5980] = 8'h00;
    mem[5981] = 8'h00;
    mem[5982] = 8'h00;
    mem[5983] = 8'h00;
    mem[5984] = 8'h00;
    mem[5985] = 8'h00;
    mem[5986] = 8'h00;
    mem[5987] = 8'h00;
    mem[5988] = 8'h00;
    mem[5989] = 8'h00;
    mem[5990] = 8'he0;
    mem[5991] = 8'hff;
    mem[5992] = 8'h03;
    mem[5993] = 8'h00;
    mem[5994] = 8'h00;
    mem[5995] = 8'hc0;
    mem[5996] = 8'hff;
    mem[5997] = 8'h3f;
    mem[5998] = 8'h00;
    mem[5999] = 8'hf0;
    mem[6000] = 8'h00;
    mem[6001] = 8'he0;
    mem[6002] = 8'h07;
    mem[6003] = 8'h3e;
    mem[6004] = 8'h00;
    mem[6005] = 8'hc0;
    mem[6006] = 8'hff;
    mem[6007] = 8'h1f;
    mem[6008] = 8'h00;
    mem[6009] = 8'h00;
    mem[6010] = 8'h00;
    mem[6011] = 8'h00;
    mem[6012] = 8'h00;
    mem[6013] = 8'h00;
    mem[6014] = 8'h00;
    mem[6015] = 8'h00;
    mem[6016] = 8'h00;
    mem[6017] = 8'h00;
    mem[6018] = 8'h00;
    mem[6019] = 8'h00;
    mem[6020] = 8'h00;
    mem[6021] = 8'h00;
    mem[6022] = 8'hc0;
    mem[6023] = 8'hff;
    mem[6024] = 8'h01;
    mem[6025] = 8'h40;
    mem[6026] = 8'h00;
    mem[6027] = 8'h00;
    mem[6028] = 8'hff;
    mem[6029] = 8'hff;
    mem[6030] = 8'h00;
    mem[6031] = 8'h00;
    mem[6032] = 8'h00;
    mem[6033] = 8'hf8;
    mem[6034] = 8'h07;
    mem[6035] = 8'h0c;
    mem[6036] = 8'h00;
    mem[6037] = 8'hf0;
    mem[6038] = 8'hff;
    mem[6039] = 8'h0f;
    mem[6040] = 8'h00;
    mem[6041] = 8'h00;
    mem[6042] = 8'h00;
    mem[6043] = 8'h00;
    mem[6044] = 8'h00;
    mem[6045] = 8'h00;
    mem[6046] = 8'h00;
    mem[6047] = 8'h00;
    mem[6048] = 8'h00;
    mem[6049] = 8'h00;
    mem[6050] = 8'h00;
    mem[6051] = 8'h00;
    mem[6052] = 8'h00;
    mem[6053] = 8'h00;
    mem[6054] = 8'h00;
    mem[6055] = 8'h7f;
    mem[6056] = 8'h00;
    mem[6057] = 8'hc0;
    mem[6058] = 8'h01;
    mem[6059] = 8'h00;
    mem[6060] = 8'hfc;
    mem[6061] = 8'hff;
    mem[6062] = 8'h03;
    mem[6063] = 8'h00;
    mem[6064] = 8'h00;
    mem[6065] = 8'hfc;
    mem[6066] = 8'h0f;
    mem[6067] = 8'h00;
    mem[6068] = 8'h00;
    mem[6069] = 8'hf8;
    mem[6070] = 8'hff;
    mem[6071] = 8'h03;
    mem[6072] = 8'h00;
    mem[6073] = 8'h00;
    mem[6074] = 8'h00;
    mem[6075] = 8'h00;
    mem[6076] = 8'h00;
    mem[6077] = 8'h00;
    mem[6078] = 8'h00;
    mem[6079] = 8'h00;
    mem[6080] = 8'h00;
    mem[6081] = 8'h00;
    mem[6082] = 8'h00;
    mem[6083] = 8'h00;
    mem[6084] = 8'h00;
    mem[6085] = 8'h00;
    mem[6086] = 8'h00;
    mem[6087] = 8'h00;
    mem[6088] = 8'h00;
    mem[6089] = 8'he0;
    mem[6090] = 8'h07;
    mem[6091] = 8'h00;
    mem[6092] = 8'hf0;
    mem[6093] = 8'hff;
    mem[6094] = 8'h0f;
    mem[6095] = 8'h00;
    mem[6096] = 8'h00;
    mem[6097] = 8'hff;
    mem[6098] = 8'h1f;
    mem[6099] = 8'h00;
    mem[6100] = 8'h00;
    mem[6101] = 8'hfe;
    mem[6102] = 8'hff;
    mem[6103] = 8'h00;
    mem[6104] = 8'h00;
    mem[6105] = 8'h00;
    mem[6106] = 8'h00;
    mem[6107] = 8'h00;
    mem[6108] = 8'h00;
    mem[6109] = 8'h00;
    mem[6110] = 8'h00;
    mem[6111] = 8'h00;
    mem[6112] = 8'h00;
    mem[6113] = 8'h00;
    mem[6114] = 8'h00;
    mem[6115] = 8'h00;
    mem[6116] = 8'h00;
    mem[6117] = 8'h00;
    mem[6118] = 8'h00;
    mem[6119] = 8'h00;
    mem[6120] = 8'h00;
    mem[6121] = 8'hf0;
    mem[6122] = 8'h0f;
    mem[6123] = 8'h00;
    mem[6124] = 8'he0;
    mem[6125] = 8'hff;
    mem[6126] = 8'h3f;
    mem[6127] = 8'h00;
    mem[6128] = 8'hc0;
    mem[6129] = 8'hff;
    mem[6130] = 8'h1f;
    mem[6131] = 8'h00;
    mem[6132] = 8'h80;
    mem[6133] = 8'hff;
    mem[6134] = 8'h7f;
    mem[6135] = 8'h00;
    mem[6136] = 8'h00;
    mem[6137] = 8'h00;
    mem[6138] = 8'h00;
    mem[6139] = 8'h00;
    mem[6140] = 8'h00;
    mem[6141] = 8'h00;
    mem[6142] = 8'h00;
    mem[6143] = 8'h00;
    mem[6144] = 8'h00;
    mem[6145] = 8'h00;
    mem[6146] = 8'h00;
    mem[6147] = 8'h00;
    mem[6148] = 8'h00;
    mem[6149] = 8'h00;
    mem[6150] = 8'h00;
    mem[6151] = 8'h00;
    mem[6152] = 8'h00;
    mem[6153] = 8'hf0;
    mem[6154] = 8'h3f;
    mem[6155] = 8'h00;
    mem[6156] = 8'h80;
    mem[6157] = 8'hff;
    mem[6158] = 8'hff;
    mem[6159] = 8'h00;
    mem[6160] = 8'hf0;
    mem[6161] = 8'hff;
    mem[6162] = 8'h3f;
    mem[6163] = 8'h00;
    mem[6164] = 8'he0;
    mem[6165] = 8'hff;
    mem[6166] = 8'h1f;
    mem[6167] = 8'h00;
    mem[6168] = 8'h00;
    mem[6169] = 8'h00;
    mem[6170] = 8'h00;
    mem[6171] = 8'h00;
    mem[6172] = 8'h00;
    mem[6173] = 8'h00;
    mem[6174] = 8'h00;
    mem[6175] = 8'h00;
    mem[6176] = 8'h00;
    mem[6177] = 8'h00;
    mem[6178] = 8'h00;
    mem[6179] = 8'h00;
    mem[6180] = 8'h00;
    mem[6181] = 8'h00;
    mem[6182] = 8'h00;
    mem[6183] = 8'h00;
    mem[6184] = 8'h00;
    mem[6185] = 8'hf8;
    mem[6186] = 8'hff;
    mem[6187] = 8'h00;
    mem[6188] = 8'h00;
    mem[6189] = 8'hfe;
    mem[6190] = 8'hff;
    mem[6191] = 8'h03;
    mem[6192] = 8'hfc;
    mem[6193] = 8'hff;
    mem[6194] = 8'h3f;
    mem[6195] = 8'h00;
    mem[6196] = 8'hf0;
    mem[6197] = 8'hff;
    mem[6198] = 8'h07;
    mem[6199] = 8'h00;
    mem[6200] = 8'h00;
    mem[6201] = 8'h00;
    mem[6202] = 8'h00;
    mem[6203] = 8'h00;
    mem[6204] = 8'h00;
    mem[6205] = 8'h00;
    mem[6206] = 8'h00;
    mem[6207] = 8'h00;
    mem[6208] = 8'h00;
    mem[6209] = 8'h00;
    mem[6210] = 8'h00;
    mem[6211] = 8'h00;
    mem[6212] = 8'h00;
    mem[6213] = 8'h00;
    mem[6214] = 8'h00;
    mem[6215] = 8'h00;
    mem[6216] = 8'h00;
    mem[6217] = 8'hf8;
    mem[6218] = 8'hff;
    mem[6219] = 8'h01;
    mem[6220] = 8'h00;
    mem[6221] = 8'hf8;
    mem[6222] = 8'hff;
    mem[6223] = 8'h8f;
    mem[6224] = 8'hff;
    mem[6225] = 8'hff;
    mem[6226] = 8'h7f;
    mem[6227] = 8'h00;
    mem[6228] = 8'hfc;
    mem[6229] = 8'hff;
    mem[6230] = 8'h03;
    mem[6231] = 8'h00;
    mem[6232] = 8'h00;
    mem[6233] = 8'h00;
    mem[6234] = 8'h00;
    mem[6235] = 8'h00;
    mem[6236] = 8'h00;
    mem[6237] = 8'h00;
    mem[6238] = 8'h00;
    mem[6239] = 8'h00;
    mem[6240] = 8'h00;
    mem[6241] = 8'h00;
    mem[6242] = 8'h00;
    mem[6243] = 8'h00;
    mem[6244] = 8'h00;
    mem[6245] = 8'h00;
    mem[6246] = 8'h00;
    mem[6247] = 8'h00;
    mem[6248] = 8'h00;
    mem[6249] = 8'hf0;
    mem[6250] = 8'hff;
    mem[6251] = 8'h07;
    mem[6252] = 8'h00;
    mem[6253] = 8'he0;
    mem[6254] = 8'hff;
    mem[6255] = 8'hff;
    mem[6256] = 8'hff;
    mem[6257] = 8'hff;
    mem[6258] = 8'hff;
    mem[6259] = 8'h00;
    mem[6260] = 8'hff;
    mem[6261] = 8'hff;
    mem[6262] = 8'h00;
    mem[6263] = 8'h00;
    mem[6264] = 8'h00;
    mem[6265] = 8'h00;
    mem[6266] = 8'h00;
    mem[6267] = 8'h00;
    mem[6268] = 8'h00;
    mem[6269] = 8'h00;
    mem[6270] = 8'h00;
    mem[6271] = 8'h00;
    mem[6272] = 8'h00;
    mem[6273] = 8'h00;
    mem[6274] = 8'h00;
    mem[6275] = 8'h00;
    mem[6276] = 8'h00;
    mem[6277] = 8'h00;
    mem[6278] = 8'h00;
    mem[6279] = 8'h00;
    mem[6280] = 8'h00;
    mem[6281] = 8'he0;
    mem[6282] = 8'hff;
    mem[6283] = 8'h1f;
    mem[6284] = 8'h00;
    mem[6285] = 8'h80;
    mem[6286] = 8'hff;
    mem[6287] = 8'hff;
    mem[6288] = 8'hff;
    mem[6289] = 8'h1f;
    mem[6290] = 8'hff;
    mem[6291] = 8'h00;
    mem[6292] = 8'hff;
    mem[6293] = 8'h3f;
    mem[6294] = 8'h00;
    mem[6295] = 8'h00;
    mem[6296] = 8'h00;
    mem[6297] = 8'h00;
    mem[6298] = 8'h00;
    mem[6299] = 8'h00;
    mem[6300] = 8'h00;
    mem[6301] = 8'h00;
    mem[6302] = 8'h00;
    mem[6303] = 8'h00;
    mem[6304] = 8'h00;
    mem[6305] = 8'h00;
    mem[6306] = 8'h00;
    mem[6307] = 8'h00;
    mem[6308] = 8'h00;
    mem[6309] = 8'h00;
    mem[6310] = 8'h00;
    mem[6311] = 8'h00;
    mem[6312] = 8'h00;
    mem[6313] = 8'h80;
    mem[6314] = 8'hff;
    mem[6315] = 8'h7f;
    mem[6316] = 8'h00;
    mem[6317] = 8'h00;
    mem[6318] = 8'hfe;
    mem[6319] = 8'hff;
    mem[6320] = 8'hff;
    mem[6321] = 8'h07;
    mem[6322] = 8'hfe;
    mem[6323] = 8'h01;
    mem[6324] = 8'hfe;
    mem[6325] = 8'h0f;
    mem[6326] = 8'h00;
    mem[6327] = 8'h00;
    mem[6328] = 8'h00;
    mem[6329] = 8'h00;
    mem[6330] = 8'h00;
    mem[6331] = 8'h00;
    mem[6332] = 8'h00;
    mem[6333] = 8'h00;
    mem[6334] = 8'h00;
    mem[6335] = 8'h00;
    mem[6336] = 8'h00;
    mem[6337] = 8'h00;
    mem[6338] = 8'h00;
    mem[6339] = 8'h00;
    mem[6340] = 8'h00;
    mem[6341] = 8'h00;
    mem[6342] = 8'h00;
    mem[6343] = 8'h00;
    mem[6344] = 8'h00;
    mem[6345] = 8'h00;
    mem[6346] = 8'hfe;
    mem[6347] = 8'hff;
    mem[6348] = 8'h01;
    mem[6349] = 8'h00;
    mem[6350] = 8'hf8;
    mem[6351] = 8'hff;
    mem[6352] = 8'hff;
    mem[6353] = 8'h01;
    mem[6354] = 8'hfe;
    mem[6355] = 8'h01;
    mem[6356] = 8'hfc;
    mem[6357] = 8'h07;
    mem[6358] = 8'h00;
    mem[6359] = 8'h00;
    mem[6360] = 8'h00;
    mem[6361] = 8'h00;
    mem[6362] = 8'h00;
    mem[6363] = 8'h00;
    mem[6364] = 8'h00;
    mem[6365] = 8'h00;
    mem[6366] = 8'h00;
    mem[6367] = 8'h00;
    mem[6368] = 8'h00;
    mem[6369] = 8'h00;
    mem[6370] = 8'h00;
    mem[6371] = 8'h00;
    mem[6372] = 8'h00;
    mem[6373] = 8'h00;
    mem[6374] = 8'h00;
    mem[6375] = 8'h00;
    mem[6376] = 8'h00;
    mem[6377] = 8'h00;
    mem[6378] = 8'hf8;
    mem[6379] = 8'hff;
    mem[6380] = 8'h03;
    mem[6381] = 8'h00;
    mem[6382] = 8'he0;
    mem[6383] = 8'hff;
    mem[6384] = 8'h7f;
    mem[6385] = 8'h00;
    mem[6386] = 8'hfc;
    mem[6387] = 8'h03;
    mem[6388] = 8'hfc;
    mem[6389] = 8'h01;
    mem[6390] = 8'h00;
    mem[6391] = 8'h00;
    mem[6392] = 8'h00;
    mem[6393] = 8'h00;
    mem[6394] = 8'h00;
    mem[6395] = 8'h00;
    mem[6396] = 8'h00;
    mem[6397] = 8'h00;
    mem[6398] = 8'h00;
    mem[6399] = 8'h00;
    mem[6400] = 8'h00;
    mem[6401] = 8'h00;
    mem[6402] = 8'h00;
    mem[6403] = 8'h00;
    mem[6404] = 8'h00;
    mem[6405] = 8'h00;
    mem[6406] = 8'h00;
    mem[6407] = 8'h00;
    mem[6408] = 8'h00;
    mem[6409] = 8'h00;
    mem[6410] = 8'hf0;
    mem[6411] = 8'hff;
    mem[6412] = 8'h0f;
    mem[6413] = 8'h00;
    mem[6414] = 8'h80;
    mem[6415] = 8'hff;
    mem[6416] = 8'h1f;
    mem[6417] = 8'h00;
    mem[6418] = 8'hfc;
    mem[6419] = 8'h07;
    mem[6420] = 8'h78;
    mem[6421] = 8'h00;
    mem[6422] = 8'h00;
    mem[6423] = 8'h00;
    mem[6424] = 8'h00;
    mem[6425] = 8'h00;
    mem[6426] = 8'h00;
    mem[6427] = 8'h00;
    mem[6428] = 8'h00;
    mem[6429] = 8'h00;
    mem[6430] = 8'h00;
    mem[6431] = 8'h00;
    mem[6432] = 8'h00;
    mem[6433] = 8'h00;
    mem[6434] = 8'h00;
    mem[6435] = 8'h00;
    mem[6436] = 8'h00;
    mem[6437] = 8'h00;
    mem[6438] = 8'h00;
    mem[6439] = 8'h00;
    mem[6440] = 8'h00;
    mem[6441] = 8'h00;
    mem[6442] = 8'hc0;
    mem[6443] = 8'hff;
    mem[6444] = 8'h3f;
    mem[6445] = 8'h00;
    mem[6446] = 8'h00;
    mem[6447] = 8'hfe;
    mem[6448] = 8'h03;
    mem[6449] = 8'h00;
    mem[6450] = 8'hf8;
    mem[6451] = 8'h07;
    mem[6452] = 8'h18;
    mem[6453] = 8'h00;
    mem[6454] = 8'h00;
    mem[6455] = 8'h00;
    mem[6456] = 8'h00;
    mem[6457] = 8'h00;
    mem[6458] = 8'h00;
    mem[6459] = 8'h00;
    mem[6460] = 8'h00;
    mem[6461] = 8'h00;
    mem[6462] = 8'h00;
    mem[6463] = 8'h00;
    mem[6464] = 8'h00;
    mem[6465] = 8'h00;
    mem[6466] = 8'h00;
    mem[6467] = 8'h00;
    mem[6468] = 8'h00;
    mem[6469] = 8'h00;
    mem[6470] = 8'h00;
    mem[6471] = 8'h00;
    mem[6472] = 8'h00;
    mem[6473] = 8'h00;
    mem[6474] = 8'h00;
    mem[6475] = 8'hff;
    mem[6476] = 8'hff;
    mem[6477] = 8'h00;
    mem[6478] = 8'h00;
    mem[6479] = 8'h70;
    mem[6480] = 8'h00;
    mem[6481] = 8'h00;
    mem[6482] = 8'hf8;
    mem[6483] = 8'h0f;
    mem[6484] = 8'h00;
    mem[6485] = 8'h00;
    mem[6486] = 8'h00;
    mem[6487] = 8'h00;
    mem[6488] = 8'h00;
    mem[6489] = 8'h00;
    mem[6490] = 8'h00;
    mem[6491] = 8'h00;
    mem[6492] = 8'h00;
    mem[6493] = 8'h00;
    mem[6494] = 8'h00;
    mem[6495] = 8'h00;
    mem[6496] = 8'h00;
    mem[6497] = 8'h00;
    mem[6498] = 8'h00;
    mem[6499] = 8'h00;
    mem[6500] = 8'h00;
    mem[6501] = 8'h00;
    mem[6502] = 8'h00;
    mem[6503] = 8'h00;
    mem[6504] = 8'h00;
    mem[6505] = 8'h00;
    mem[6506] = 8'h00;
    mem[6507] = 8'hfc;
    mem[6508] = 8'hff;
    mem[6509] = 8'h03;
    mem[6510] = 8'h00;
    mem[6511] = 8'h00;
    mem[6512] = 8'h00;
    mem[6513] = 8'h00;
    mem[6514] = 8'hfc;
    mem[6515] = 8'h0f;
    mem[6516] = 8'h00;
    mem[6517] = 8'h00;
    mem[6518] = 8'h00;
    mem[6519] = 8'h00;
    mem[6520] = 8'h00;
    mem[6521] = 8'h00;
    mem[6522] = 8'h00;
    mem[6523] = 8'h00;
    mem[6524] = 8'h00;
    mem[6525] = 8'h00;
    mem[6526] = 8'h00;
    mem[6527] = 8'h00;
    mem[6528] = 8'h00;
    mem[6529] = 8'h00;
    mem[6530] = 8'h00;
    mem[6531] = 8'h00;
    mem[6532] = 8'h00;
    mem[6533] = 8'h00;
    mem[6534] = 8'h00;
    mem[6535] = 8'h00;
    mem[6536] = 8'h00;
    mem[6537] = 8'h00;
    mem[6538] = 8'h00;
    mem[6539] = 8'hf0;
    mem[6540] = 8'hff;
    mem[6541] = 8'h0f;
    mem[6542] = 8'h00;
    mem[6543] = 8'h00;
    mem[6544] = 8'h00;
    mem[6545] = 8'h00;
    mem[6546] = 8'hff;
    mem[6547] = 8'h1f;
    mem[6548] = 8'h00;
    mem[6549] = 8'h00;
    mem[6550] = 8'h00;
    mem[6551] = 8'h00;
    mem[6552] = 8'h00;
    mem[6553] = 8'h00;
    mem[6554] = 8'h00;
    mem[6555] = 8'h00;
    mem[6556] = 8'h00;
    mem[6557] = 8'h00;
    mem[6558] = 8'h00;
    mem[6559] = 8'h00;
    mem[6560] = 8'h00;
    mem[6561] = 8'h00;
    mem[6562] = 8'h00;
    mem[6563] = 8'h00;
    mem[6564] = 8'h00;
    mem[6565] = 8'h00;
    mem[6566] = 8'h00;
    mem[6567] = 8'h00;
    mem[6568] = 8'h00;
    mem[6569] = 8'h00;
    mem[6570] = 8'h00;
    mem[6571] = 8'he0;
    mem[6572] = 8'hff;
    mem[6573] = 8'h1f;
    mem[6574] = 8'h00;
    mem[6575] = 8'h00;
    mem[6576] = 8'h00;
    mem[6577] = 8'hc0;
    mem[6578] = 8'hff;
    mem[6579] = 8'h1f;
    mem[6580] = 8'h00;
    mem[6581] = 8'h00;
    mem[6582] = 8'h00;
    mem[6583] = 8'h00;
    mem[6584] = 8'h00;
    mem[6585] = 8'h00;
    mem[6586] = 8'h00;
    mem[6587] = 8'h00;
    mem[6588] = 8'h00;
    mem[6589] = 8'h00;
    mem[6590] = 8'h00;
    mem[6591] = 8'h00;
    mem[6592] = 8'h00;
    mem[6593] = 8'h00;
    mem[6594] = 8'h00;
    mem[6595] = 8'h00;
    mem[6596] = 8'h00;
    mem[6597] = 8'h00;
    mem[6598] = 8'h00;
    mem[6599] = 8'h00;
    mem[6600] = 8'h00;
    mem[6601] = 8'h00;
    mem[6602] = 8'h00;
    mem[6603] = 8'h80;
    mem[6604] = 8'hff;
    mem[6605] = 8'h7f;
    mem[6606] = 8'h00;
    mem[6607] = 8'h00;
    mem[6608] = 8'h00;
    mem[6609] = 8'hf0;
    mem[6610] = 8'hff;
    mem[6611] = 8'h1f;
    mem[6612] = 8'h00;
    mem[6613] = 8'h00;
    mem[6614] = 8'h00;
    mem[6615] = 8'h00;
    mem[6616] = 8'h00;
    mem[6617] = 8'h00;
    mem[6618] = 8'h00;
    mem[6619] = 8'h00;
    mem[6620] = 8'h00;
    mem[6621] = 8'h00;
    mem[6622] = 8'h00;
    mem[6623] = 8'h00;
    mem[6624] = 8'h00;
    mem[6625] = 8'h00;
    mem[6626] = 8'h00;
    mem[6627] = 8'h00;
    mem[6628] = 8'h00;
    mem[6629] = 8'h00;
    mem[6630] = 8'h00;
    mem[6631] = 8'h00;
    mem[6632] = 8'h00;
    mem[6633] = 8'h00;
    mem[6634] = 8'h00;
    mem[6635] = 8'h00;
    mem[6636] = 8'hfe;
    mem[6637] = 8'hff;
    mem[6638] = 8'h01;
    mem[6639] = 8'h00;
    mem[6640] = 8'h00;
    mem[6641] = 8'hfc;
    mem[6642] = 8'hff;
    mem[6643] = 8'h07;
    mem[6644] = 8'h00;
    mem[6645] = 8'h00;
    mem[6646] = 8'h00;
    mem[6647] = 8'h00;
    mem[6648] = 8'h00;
    mem[6649] = 8'h00;
    mem[6650] = 8'h00;
    mem[6651] = 8'h00;
    mem[6652] = 8'h00;
    mem[6653] = 8'h00;
    mem[6654] = 8'h00;
    mem[6655] = 8'h00;
    mem[6656] = 8'h00;
    mem[6657] = 8'h00;
    mem[6658] = 8'h00;
    mem[6659] = 8'h00;
    mem[6660] = 8'h00;
    mem[6661] = 8'h00;
    mem[6662] = 8'h00;
    mem[6663] = 8'h00;
    mem[6664] = 8'h00;
    mem[6665] = 8'h00;
    mem[6666] = 8'h00;
    mem[6667] = 8'h00;
    mem[6668] = 8'hf8;
    mem[6669] = 8'hff;
    mem[6670] = 8'h07;
    mem[6671] = 8'h00;
    mem[6672] = 8'h00;
    mem[6673] = 8'hff;
    mem[6674] = 8'hff;
    mem[6675] = 8'h01;
    mem[6676] = 8'h00;
    mem[6677] = 8'h00;
    mem[6678] = 8'h00;
    mem[6679] = 8'h00;
    mem[6680] = 8'h00;
    mem[6681] = 8'h00;
    mem[6682] = 8'h00;
    mem[6683] = 8'h00;
    mem[6684] = 8'h00;
    mem[6685] = 8'h00;
    mem[6686] = 8'h00;
    mem[6687] = 8'h00;
    mem[6688] = 8'h00;
    mem[6689] = 8'h00;
    mem[6690] = 8'h00;
    mem[6691] = 8'h00;
    mem[6692] = 8'h00;
    mem[6693] = 8'h00;
    mem[6694] = 8'h00;
    mem[6695] = 8'h00;
    mem[6696] = 8'h00;
    mem[6697] = 8'h00;
    mem[6698] = 8'h00;
    mem[6699] = 8'h00;
    mem[6700] = 8'he0;
    mem[6701] = 8'hff;
    mem[6702] = 8'h1f;
    mem[6703] = 8'h00;
    mem[6704] = 8'hc0;
    mem[6705] = 8'hff;
    mem[6706] = 8'h7f;
    mem[6707] = 8'h00;
    mem[6708] = 8'h00;
    mem[6709] = 8'h00;
    mem[6710] = 8'h00;
    mem[6711] = 8'h00;
    mem[6712] = 8'h00;
    mem[6713] = 8'h00;
    mem[6714] = 8'h00;
    mem[6715] = 8'h00;
    mem[6716] = 8'h00;
    mem[6717] = 8'h00;
    mem[6718] = 8'h00;
    mem[6719] = 8'h00;
    mem[6720] = 8'h00;
    mem[6721] = 8'h00;
    mem[6722] = 8'h00;
    mem[6723] = 8'h00;
    mem[6724] = 8'h00;
    mem[6725] = 8'h00;
    mem[6726] = 8'h00;
    mem[6727] = 8'h00;
    mem[6728] = 8'h00;
    mem[6729] = 8'h00;
    mem[6730] = 8'h00;
    mem[6731] = 8'h00;
    mem[6732] = 8'h80;
    mem[6733] = 8'hff;
    mem[6734] = 8'h7f;
    mem[6735] = 8'h00;
    mem[6736] = 8'hf0;
    mem[6737] = 8'hff;
    mem[6738] = 8'h1f;
    mem[6739] = 8'h00;
    mem[6740] = 8'h00;
    mem[6741] = 8'h00;
    mem[6742] = 8'h00;
    mem[6743] = 8'h00;
    mem[6744] = 8'h00;
    mem[6745] = 8'h00;
    mem[6746] = 8'h00;
    mem[6747] = 8'h00;
    mem[6748] = 8'h00;
    mem[6749] = 8'h00;
    mem[6750] = 8'h00;
    mem[6751] = 8'h00;
    mem[6752] = 8'h00;
    mem[6753] = 8'h00;
    mem[6754] = 8'h00;
    mem[6755] = 8'h00;
    mem[6756] = 8'h00;
    mem[6757] = 8'h00;
    mem[6758] = 8'h00;
    mem[6759] = 8'h00;
    mem[6760] = 8'h00;
    mem[6761] = 8'h00;
    mem[6762] = 8'h00;
    mem[6763] = 8'h00;
    mem[6764] = 8'h00;
    mem[6765] = 8'hfe;
    mem[6766] = 8'hff;
    mem[6767] = 8'h01;
    mem[6768] = 8'hfc;
    mem[6769] = 8'hff;
    mem[6770] = 8'h07;
    mem[6771] = 8'h00;
    mem[6772] = 8'h00;
    mem[6773] = 8'h00;
    mem[6774] = 8'h00;
    mem[6775] = 8'h00;
    mem[6776] = 8'h00;
    mem[6777] = 8'h00;
    mem[6778] = 8'h00;
    mem[6779] = 8'h00;
    mem[6780] = 8'h00;
    mem[6781] = 8'h00;
    mem[6782] = 8'h00;
    mem[6783] = 8'h00;
    mem[6784] = 8'h00;
    mem[6785] = 8'h00;
    mem[6786] = 8'h00;
    mem[6787] = 8'h00;
    mem[6788] = 8'h00;
    mem[6789] = 8'h00;
    mem[6790] = 8'h00;
    mem[6791] = 8'h00;
    mem[6792] = 8'h00;
    mem[6793] = 8'h00;
    mem[6794] = 8'h00;
    mem[6795] = 8'h00;
    mem[6796] = 8'h00;
    mem[6797] = 8'hfc;
    mem[6798] = 8'hff;
    mem[6799] = 8'h0f;
    mem[6800] = 8'hff;
    mem[6801] = 8'hff;
    mem[6802] = 8'h01;
    mem[6803] = 8'h00;
    mem[6804] = 8'h00;
    mem[6805] = 8'h00;
    mem[6806] = 8'h00;
    mem[6807] = 8'h00;
    mem[6808] = 8'h00;
    mem[6809] = 8'h00;
    mem[6810] = 8'h00;
    mem[6811] = 8'h00;
    mem[6812] = 8'h00;
    mem[6813] = 8'h00;
    mem[6814] = 8'h00;
    mem[6815] = 8'h00;
    mem[6816] = 8'h00;
    mem[6817] = 8'h00;
    mem[6818] = 8'h00;
    mem[6819] = 8'h00;
    mem[6820] = 8'h00;
    mem[6821] = 8'h00;
    mem[6822] = 8'h00;
    mem[6823] = 8'h00;
    mem[6824] = 8'h00;
    mem[6825] = 8'h00;
    mem[6826] = 8'h00;
    mem[6827] = 8'h00;
    mem[6828] = 8'h00;
    mem[6829] = 8'hf0;
    mem[6830] = 8'hff;
    mem[6831] = 8'hff;
    mem[6832] = 8'hff;
    mem[6833] = 8'h7f;
    mem[6834] = 8'h00;
    mem[6835] = 8'h00;
    mem[6836] = 8'h00;
    mem[6837] = 8'h00;
    mem[6838] = 8'h00;
    mem[6839] = 8'h00;
    mem[6840] = 8'h00;
    mem[6841] = 8'h00;
    mem[6842] = 8'h00;
    mem[6843] = 8'h00;
    mem[6844] = 8'h00;
    mem[6845] = 8'h00;
    mem[6846] = 8'h00;
    mem[6847] = 8'h00;
    mem[6848] = 8'h00;
    mem[6849] = 8'h00;
    mem[6850] = 8'h00;
    mem[6851] = 8'h00;
    mem[6852] = 8'h00;
    mem[6853] = 8'h00;
    mem[6854] = 8'h00;
    mem[6855] = 8'h00;
    mem[6856] = 8'h00;
    mem[6857] = 8'h00;
    mem[6858] = 8'h00;
    mem[6859] = 8'h00;
    mem[6860] = 8'h00;
    mem[6861] = 8'hc0;
    mem[6862] = 8'hff;
    mem[6863] = 8'hff;
    mem[6864] = 8'hff;
    mem[6865] = 8'h1f;
    mem[6866] = 8'h00;
    mem[6867] = 8'h00;
    mem[6868] = 8'h00;
    mem[6869] = 8'h00;
    mem[6870] = 8'h00;
    mem[6871] = 8'h00;
    mem[6872] = 8'h00;
    mem[6873] = 8'h00;
    mem[6874] = 8'h00;
    mem[6875] = 8'h00;
    mem[6876] = 8'h00;
    mem[6877] = 8'h00;
    mem[6878] = 8'h00;
    mem[6879] = 8'h00;
    mem[6880] = 8'h00;
    mem[6881] = 8'h00;
    mem[6882] = 8'h00;
    mem[6883] = 8'h00;
    mem[6884] = 8'h00;
    mem[6885] = 8'h00;
    mem[6886] = 8'h00;
    mem[6887] = 8'h00;
    mem[6888] = 8'h00;
    mem[6889] = 8'h00;
    mem[6890] = 8'h00;
    mem[6891] = 8'h00;
    mem[6892] = 8'h00;
    mem[6893] = 8'h00;
    mem[6894] = 8'hff;
    mem[6895] = 8'hff;
    mem[6896] = 8'hff;
    mem[6897] = 8'h07;
    mem[6898] = 8'h00;
    mem[6899] = 8'h00;
    mem[6900] = 8'h00;
    mem[6901] = 8'h00;
    mem[6902] = 8'h00;
    mem[6903] = 8'h00;
    mem[6904] = 8'h00;
    mem[6905] = 8'h00;
    mem[6906] = 8'h00;
    mem[6907] = 8'h00;
    mem[6908] = 8'h00;
    mem[6909] = 8'h00;
    mem[6910] = 8'h00;
    mem[6911] = 8'h00;
    mem[6912] = 8'h00;
    mem[6913] = 8'h00;
    mem[6914] = 8'h00;
    mem[6915] = 8'h00;
    mem[6916] = 8'h00;
    mem[6917] = 8'h00;
    mem[6918] = 8'h00;
    mem[6919] = 8'h00;
    mem[6920] = 8'h00;
    mem[6921] = 8'h00;
    mem[6922] = 8'h00;
    mem[6923] = 8'h00;
    mem[6924] = 8'h00;
    mem[6925] = 8'h00;
    mem[6926] = 8'hf8;
    mem[6927] = 8'hff;
    mem[6928] = 8'hff;
    mem[6929] = 8'h01;
    mem[6930] = 8'h00;
    mem[6931] = 8'h00;
    mem[6932] = 8'h00;
    mem[6933] = 8'h00;
    mem[6934] = 8'h00;
    mem[6935] = 8'h00;
    mem[6936] = 8'h00;
    mem[6937] = 8'h00;
    mem[6938] = 8'h00;
    mem[6939] = 8'h00;
    mem[6940] = 8'h00;
    mem[6941] = 8'h00;
    mem[6942] = 8'h00;
    mem[6943] = 8'h00;
    mem[6944] = 8'h00;
    mem[6945] = 8'h00;
    mem[6946] = 8'h00;
    mem[6947] = 8'h00;
    mem[6948] = 8'h00;
    mem[6949] = 8'h00;
    mem[6950] = 8'h00;
    mem[6951] = 8'h00;
    mem[6952] = 8'h00;
    mem[6953] = 8'h00;
    mem[6954] = 8'h00;
    mem[6955] = 8'h00;
    mem[6956] = 8'h00;
    mem[6957] = 8'h00;
    mem[6958] = 8'he0;
    mem[6959] = 8'hff;
    mem[6960] = 8'h7f;
    mem[6961] = 8'h00;
    mem[6962] = 8'h00;
    mem[6963] = 8'h00;
    mem[6964] = 8'h00;
    mem[6965] = 8'h00;
    mem[6966] = 8'h00;
    mem[6967] = 8'h00;
    mem[6968] = 8'h00;
    mem[6969] = 8'h00;
    mem[6970] = 8'h00;
    mem[6971] = 8'h00;
    mem[6972] = 8'h00;
    mem[6973] = 8'h00;
    mem[6974] = 8'h00;
    mem[6975] = 8'h00;
    mem[6976] = 8'h00;
    mem[6977] = 8'h00;
    mem[6978] = 8'h00;
    mem[6979] = 8'h00;
    mem[6980] = 8'h00;
    mem[6981] = 8'h00;
    mem[6982] = 8'h00;
    mem[6983] = 8'h00;
    mem[6984] = 8'h00;
    mem[6985] = 8'h00;
    mem[6986] = 8'h00;
    mem[6987] = 8'h00;
    mem[6988] = 8'h00;
    mem[6989] = 8'h00;
    mem[6990] = 8'h80;
    mem[6991] = 8'hff;
    mem[6992] = 8'h1f;
    mem[6993] = 8'h00;
    mem[6994] = 8'h00;
    mem[6995] = 8'h00;
    mem[6996] = 8'h00;
    mem[6997] = 8'h00;
    mem[6998] = 8'h00;
    mem[6999] = 8'h00;
    mem[7000] = 8'h00;
    mem[7001] = 8'h00;
    mem[7002] = 8'h00;
    mem[7003] = 8'h00;
    mem[7004] = 8'h00;
    mem[7005] = 8'h00;
    mem[7006] = 8'h00;
    mem[7007] = 8'h00;
    mem[7008] = 8'h00;
    mem[7009] = 8'h00;
    mem[7010] = 8'h00;
    mem[7011] = 8'h00;
    mem[7012] = 8'h00;
    mem[7013] = 8'h00;
    mem[7014] = 8'h00;
    mem[7015] = 8'h00;
    mem[7016] = 8'h00;
    mem[7017] = 8'h00;
    mem[7018] = 8'h00;
    mem[7019] = 8'h00;
    mem[7020] = 8'h00;
    mem[7021] = 8'h00;
    mem[7022] = 8'h00;
    mem[7023] = 8'hfe;
    mem[7024] = 8'h03;
    mem[7025] = 8'h00;
    mem[7026] = 8'h00;
    mem[7027] = 8'h00;
    mem[7028] = 8'h00;
    mem[7029] = 8'h00;
    mem[7030] = 8'h00;
    mem[7031] = 8'h00;
    mem[7032] = 8'h00;
    mem[7033] = 8'h00;
    mem[7034] = 8'h00;
    mem[7035] = 8'h00;
    mem[7036] = 8'h00;
    mem[7037] = 8'h00;
    mem[7038] = 8'h00;
    mem[7039] = 8'h00;
    mem[7040] = 8'h00;
    mem[7041] = 8'h00;
    mem[7042] = 8'h00;
    mem[7043] = 8'h00;
    mem[7044] = 8'h00;
    mem[7045] = 8'h00;
    mem[7046] = 8'h00;
    mem[7047] = 8'h00;
    mem[7048] = 8'h00;
    mem[7049] = 8'h00;
    mem[7050] = 8'h00;
    mem[7051] = 8'h00;
    mem[7052] = 8'h00;
    mem[7053] = 8'h00;
    mem[7054] = 8'h00;
    mem[7055] = 8'hf0;
    mem[7056] = 8'h00;
    mem[7057] = 8'h00;
    mem[7058] = 8'h00;
    mem[7059] = 8'h00;
    mem[7060] = 8'h00;
    mem[7061] = 8'h00;
    mem[7062] = 8'h00;
    mem[7063] = 8'h00;
    mem[7064] = 8'h00;
    mem[7065] = 8'h00;
    mem[7066] = 8'h00;
    mem[7067] = 8'h00;
    mem[7068] = 8'h00;
    mem[7069] = 8'h00;
    mem[7070] = 8'h00;
    mem[7071] = 8'h00;
    mem[7072] = 8'h00;
    mem[7073] = 8'h00;
    mem[7074] = 8'h00;
    mem[7075] = 8'h00;
    mem[7076] = 8'h00;
    mem[7077] = 8'h00;
    mem[7078] = 8'h00;
    mem[7079] = 8'h00;
    mem[7080] = 8'h00;
    mem[7081] = 8'h00;
    mem[7082] = 8'h00;
    mem[7083] = 8'h00;
    mem[7084] = 8'h00;
    mem[7085] = 8'h00;
    mem[7086] = 8'h00;
    mem[7087] = 8'h00;
    mem[7088] = 8'h00;
    mem[7089] = 8'h00;
    mem[7090] = 8'h00;
    mem[7091] = 8'h00;
    mem[7092] = 8'h00;
    mem[7093] = 8'h00;
    mem[7094] = 8'h00;
    mem[7095] = 8'h00;
    mem[7096] = 8'h00;
    mem[7097] = 8'h00;
    mem[7098] = 8'h00;
    mem[7099] = 8'h00;
    mem[7100] = 8'h00;
    mem[7101] = 8'h00;
    mem[7102] = 8'h00;
    mem[7103] = 8'h00;
    mem[7104] = 8'h00;
    mem[7105] = 8'h00;
    mem[7106] = 8'h00;
    mem[7107] = 8'h00;
    mem[7108] = 8'h00;
    mem[7109] = 8'h00;
    mem[7110] = 8'h00;
    mem[7111] = 8'h00;
    mem[7112] = 8'h00;
    mem[7113] = 8'h00;
    mem[7114] = 8'h00;
    mem[7115] = 8'h00;
    mem[7116] = 8'h00;
    mem[7117] = 8'h00;
    mem[7118] = 8'h00;
    mem[7119] = 8'h00;
    mem[7120] = 8'h00;
    mem[7121] = 8'h00;
    mem[7122] = 8'h00;
    mem[7123] = 8'h00;
    mem[7124] = 8'h00;
    mem[7125] = 8'h00;
    mem[7126] = 8'h00;
    mem[7127] = 8'h00;
    mem[7128] = 8'h00;
    mem[7129] = 8'h00;
    mem[7130] = 8'h00;
    mem[7131] = 8'h00;
    mem[7132] = 8'h00;
    mem[7133] = 8'h00;
    mem[7134] = 8'h00;
    mem[7135] = 8'h00;
    mem[7136] = 8'h00;
    mem[7137] = 8'h00;
    mem[7138] = 8'h00;
    mem[7139] = 8'h00;
    mem[7140] = 8'h00;
    mem[7141] = 8'h00;
    mem[7142] = 8'h00;
    mem[7143] = 8'h00;
    mem[7144] = 8'h00;
    mem[7145] = 8'h00;
    mem[7146] = 8'h00;
    mem[7147] = 8'he0;
    mem[7148] = 8'h00;
    mem[7149] = 8'h00;
    mem[7150] = 8'h00;
    mem[7151] = 8'h00;
    mem[7152] = 8'h00;
    mem[7153] = 8'h00;
    mem[7154] = 8'h07;
    mem[7155] = 8'h00;
    mem[7156] = 8'h00;
    mem[7157] = 8'h00;
    mem[7158] = 8'h00;
    mem[7159] = 8'h0f;
    mem[7160] = 8'h00;
    mem[7161] = 8'h0f;
    mem[7162] = 8'h00;
    mem[7163] = 8'h00;
    mem[7164] = 8'h00;
    mem[7165] = 8'h00;
    mem[7166] = 8'h00;
    mem[7167] = 8'h00;
    mem[7168] = 8'h00;
    mem[7169] = 8'h00;
    mem[7170] = 8'h00;
    mem[7171] = 8'h00;
    mem[7172] = 8'h00;
    mem[7173] = 8'hfe;
    mem[7174] = 8'h9f;
    mem[7175] = 8'hff;
    mem[7176] = 8'h03;
    mem[7177] = 8'h07;
    mem[7178] = 8'h0e;
    mem[7179] = 8'hfc;
    mem[7180] = 8'h07;
    mem[7181] = 8'hf0;
    mem[7182] = 8'he0;
    mem[7183] = 8'hff;
    mem[7184] = 8'h73;
    mem[7185] = 8'he0;
    mem[7186] = 8'h3f;
    mem[7187] = 8'hf0;
    mem[7188] = 8'hc0;
    mem[7189] = 8'h01;
    mem[7190] = 8'he0;
    mem[7191] = 8'h3f;
    mem[7192] = 8'hc0;
    mem[7193] = 8'h7f;
    mem[7194] = 8'h00;
    mem[7195] = 8'h00;
    mem[7196] = 8'h00;
    mem[7197] = 8'h00;
    mem[7198] = 8'h00;
    mem[7199] = 8'h00;
    mem[7200] = 8'h00;
    mem[7201] = 8'h00;
    mem[7202] = 8'h00;
    mem[7203] = 8'h00;
    mem[7204] = 8'h00;
    mem[7205] = 8'hfe;
    mem[7206] = 8'h9f;
    mem[7207] = 8'hff;
    mem[7208] = 8'h07;
    mem[7209] = 8'h07;
    mem[7210] = 8'h0e;
    mem[7211] = 8'hfe;
    mem[7212] = 8'h0f;
    mem[7213] = 8'hf8;
    mem[7214] = 8'he0;
    mem[7215] = 8'hff;
    mem[7216] = 8'h73;
    mem[7217] = 8'hf0;
    mem[7218] = 8'h7f;
    mem[7219] = 8'hf0;
    mem[7220] = 8'hc0;
    mem[7221] = 8'h01;
    mem[7222] = 8'hf0;
    mem[7223] = 8'h7f;
    mem[7224] = 8'he0;
    mem[7225] = 8'hff;
    mem[7226] = 8'h00;
    mem[7227] = 8'h00;
    mem[7228] = 8'h00;
    mem[7229] = 8'h00;
    mem[7230] = 8'h00;
    mem[7231] = 8'h00;
    mem[7232] = 8'h00;
    mem[7233] = 8'h00;
    mem[7234] = 8'h00;
    mem[7235] = 8'h00;
    mem[7236] = 8'h00;
    mem[7237] = 8'hfe;
    mem[7238] = 8'h9f;
    mem[7239] = 8'hff;
    mem[7240] = 8'h0f;
    mem[7241] = 8'h07;
    mem[7242] = 8'h0e;
    mem[7243] = 8'h1f;
    mem[7244] = 8'h1f;
    mem[7245] = 8'hf8;
    mem[7246] = 8'he1;
    mem[7247] = 8'hff;
    mem[7248] = 8'h73;
    mem[7249] = 8'hf8;
    mem[7250] = 8'hf8;
    mem[7251] = 8'hf0;
    mem[7252] = 8'hc1;
    mem[7253] = 8'h01;
    mem[7254] = 8'hf8;
    mem[7255] = 8'hf8;
    mem[7256] = 8'hf0;
    mem[7257] = 8'hf1;
    mem[7258] = 8'h01;
    mem[7259] = 8'h00;
    mem[7260] = 8'h00;
    mem[7261] = 8'h00;
    mem[7262] = 8'h00;
    mem[7263] = 8'h00;
    mem[7264] = 8'h00;
    mem[7265] = 8'h00;
    mem[7266] = 8'h00;
    mem[7267] = 8'h00;
    mem[7268] = 8'h00;
    mem[7269] = 8'h0e;
    mem[7270] = 8'h80;
    mem[7271] = 8'h07;
    mem[7272] = 8'h0f;
    mem[7273] = 8'h07;
    mem[7274] = 8'h0e;
    mem[7275] = 8'h07;
    mem[7276] = 8'h1c;
    mem[7277] = 8'hf8;
    mem[7278] = 8'h01;
    mem[7279] = 8'h1c;
    mem[7280] = 8'h70;
    mem[7281] = 8'h38;
    mem[7282] = 8'he0;
    mem[7283] = 8'hf0;
    mem[7284] = 8'hc3;
    mem[7285] = 8'h01;
    mem[7286] = 8'h78;
    mem[7287] = 8'he0;
    mem[7288] = 8'h78;
    mem[7289] = 8'hc0;
    mem[7290] = 8'h01;
    mem[7291] = 8'h00;
    mem[7292] = 8'h00;
    mem[7293] = 8'h00;
    mem[7294] = 8'h00;
    mem[7295] = 8'h00;
    mem[7296] = 8'h00;
    mem[7297] = 8'h00;
    mem[7298] = 8'h00;
    mem[7299] = 8'h00;
    mem[7300] = 8'h00;
    mem[7301] = 8'h0e;
    mem[7302] = 8'h80;
    mem[7303] = 8'h07;
    mem[7304] = 8'h1e;
    mem[7305] = 8'h07;
    mem[7306] = 8'h8e;
    mem[7307] = 8'h07;
    mem[7308] = 8'h1c;
    mem[7309] = 8'hdc;
    mem[7310] = 8'h03;
    mem[7311] = 8'h1c;
    mem[7312] = 8'h70;
    mem[7313] = 8'h3c;
    mem[7314] = 8'he0;
    mem[7315] = 8'hf1;
    mem[7316] = 8'hc3;
    mem[7317] = 8'h01;
    mem[7318] = 8'h3c;
    mem[7319] = 8'he0;
    mem[7320] = 8'h38;
    mem[7321] = 8'hc0;
    mem[7322] = 8'h03;
    mem[7323] = 8'h00;
    mem[7324] = 8'h00;
    mem[7325] = 8'h00;
    mem[7326] = 8'h00;
    mem[7327] = 8'h00;
    mem[7328] = 8'h00;
    mem[7329] = 8'h00;
    mem[7330] = 8'h00;
    mem[7331] = 8'h00;
    mem[7332] = 8'h00;
    mem[7333] = 8'h0e;
    mem[7334] = 8'h80;
    mem[7335] = 8'h07;
    mem[7336] = 8'h1e;
    mem[7337] = 8'h07;
    mem[7338] = 8'h8e;
    mem[7339] = 8'h03;
    mem[7340] = 8'h00;
    mem[7341] = 8'h9c;
    mem[7342] = 8'h03;
    mem[7343] = 8'h1c;
    mem[7344] = 8'h70;
    mem[7345] = 8'h1c;
    mem[7346] = 8'hc0;
    mem[7347] = 8'h71;
    mem[7348] = 8'hc7;
    mem[7349] = 8'h01;
    mem[7350] = 8'h3c;
    mem[7351] = 8'h00;
    mem[7352] = 8'h38;
    mem[7353] = 8'hc0;
    mem[7354] = 8'h03;
    mem[7355] = 8'h00;
    mem[7356] = 8'h00;
    mem[7357] = 8'h00;
    mem[7358] = 8'h00;
    mem[7359] = 8'h00;
    mem[7360] = 8'h00;
    mem[7361] = 8'h00;
    mem[7362] = 8'h00;
    mem[7363] = 8'h00;
    mem[7364] = 8'h00;
    mem[7365] = 8'hfe;
    mem[7366] = 8'h8f;
    mem[7367] = 8'h07;
    mem[7368] = 8'h1c;
    mem[7369] = 8'h07;
    mem[7370] = 8'h8e;
    mem[7371] = 8'h03;
    mem[7372] = 8'h00;
    mem[7373] = 8'h9c;
    mem[7374] = 8'h03;
    mem[7375] = 8'h1c;
    mem[7376] = 8'h70;
    mem[7377] = 8'h1c;
    mem[7378] = 8'hc0;
    mem[7379] = 8'h71;
    mem[7380] = 8'hc7;
    mem[7381] = 8'h01;
    mem[7382] = 8'h1c;
    mem[7383] = 8'h00;
    mem[7384] = 8'h38;
    mem[7385] = 8'h80;
    mem[7386] = 8'h03;
    mem[7387] = 8'h00;
    mem[7388] = 8'h00;
    mem[7389] = 8'h00;
    mem[7390] = 8'h00;
    mem[7391] = 8'h00;
    mem[7392] = 8'h00;
    mem[7393] = 8'h00;
    mem[7394] = 8'h00;
    mem[7395] = 8'h00;
    mem[7396] = 8'h00;
    mem[7397] = 8'hfe;
    mem[7398] = 8'h8f;
    mem[7399] = 8'h07;
    mem[7400] = 8'h1c;
    mem[7401] = 8'h07;
    mem[7402] = 8'h8e;
    mem[7403] = 8'h03;
    mem[7404] = 8'h00;
    mem[7405] = 8'h8e;
    mem[7406] = 8'h07;
    mem[7407] = 8'h1c;
    mem[7408] = 8'h70;
    mem[7409] = 8'h1c;
    mem[7410] = 8'hc0;
    mem[7411] = 8'h71;
    mem[7412] = 8'hce;
    mem[7413] = 8'h01;
    mem[7414] = 8'h1c;
    mem[7415] = 8'h00;
    mem[7416] = 8'h3c;
    mem[7417] = 8'h80;
    mem[7418] = 8'h03;
    mem[7419] = 8'h00;
    mem[7420] = 8'h00;
    mem[7421] = 8'h00;
    mem[7422] = 8'h00;
    mem[7423] = 8'h00;
    mem[7424] = 8'h00;
    mem[7425] = 8'h00;
    mem[7426] = 8'h00;
    mem[7427] = 8'h00;
    mem[7428] = 8'h00;
    mem[7429] = 8'hfe;
    mem[7430] = 8'h8f;
    mem[7431] = 8'h07;
    mem[7432] = 8'h1c;
    mem[7433] = 8'h07;
    mem[7434] = 8'h8e;
    mem[7435] = 8'h03;
    mem[7436] = 8'h00;
    mem[7437] = 8'h0e;
    mem[7438] = 8'h07;
    mem[7439] = 8'h1c;
    mem[7440] = 8'h70;
    mem[7441] = 8'h1c;
    mem[7442] = 8'hc0;
    mem[7443] = 8'h71;
    mem[7444] = 8'hde;
    mem[7445] = 8'h01;
    mem[7446] = 8'h1c;
    mem[7447] = 8'h00;
    mem[7448] = 8'h38;
    mem[7449] = 8'h80;
    mem[7450] = 8'h03;
    mem[7451] = 8'h00;
    mem[7452] = 8'h00;
    mem[7453] = 8'h00;
    mem[7454] = 8'h00;
    mem[7455] = 8'h00;
    mem[7456] = 8'h00;
    mem[7457] = 8'h00;
    mem[7458] = 8'h00;
    mem[7459] = 8'h00;
    mem[7460] = 8'h00;
    mem[7461] = 8'h0e;
    mem[7462] = 8'h80;
    mem[7463] = 8'h07;
    mem[7464] = 8'h1e;
    mem[7465] = 8'h07;
    mem[7466] = 8'h8e;
    mem[7467] = 8'h03;
    mem[7468] = 8'h00;
    mem[7469] = 8'h0e;
    mem[7470] = 8'h07;
    mem[7471] = 8'h1c;
    mem[7472] = 8'h70;
    mem[7473] = 8'h1c;
    mem[7474] = 8'hc0;
    mem[7475] = 8'h71;
    mem[7476] = 8'hdc;
    mem[7477] = 8'h01;
    mem[7478] = 8'h1c;
    mem[7479] = 8'h00;
    mem[7480] = 8'h38;
    mem[7481] = 8'h80;
    mem[7482] = 8'h03;
    mem[7483] = 8'h00;
    mem[7484] = 8'h00;
    mem[7485] = 8'h00;
    mem[7486] = 8'h00;
    mem[7487] = 8'h00;
    mem[7488] = 8'h00;
    mem[7489] = 8'h00;
    mem[7490] = 8'h00;
    mem[7491] = 8'h00;
    mem[7492] = 8'h00;
    mem[7493] = 8'h0e;
    mem[7494] = 8'h80;
    mem[7495] = 8'h07;
    mem[7496] = 8'h1e;
    mem[7497] = 8'h07;
    mem[7498] = 8'h8e;
    mem[7499] = 8'h07;
    mem[7500] = 8'h1c;
    mem[7501] = 8'hff;
    mem[7502] = 8'h0f;
    mem[7503] = 8'h1c;
    mem[7504] = 8'h70;
    mem[7505] = 8'h3c;
    mem[7506] = 8'hc0;
    mem[7507] = 8'h71;
    mem[7508] = 8'hf8;
    mem[7509] = 8'h01;
    mem[7510] = 8'h3c;
    mem[7511] = 8'he0;
    mem[7512] = 8'h39;
    mem[7513] = 8'hc0;
    mem[7514] = 8'h03;
    mem[7515] = 8'h00;
    mem[7516] = 8'h00;
    mem[7517] = 8'h00;
    mem[7518] = 8'h00;
    mem[7519] = 8'h00;
    mem[7520] = 8'h00;
    mem[7521] = 8'h00;
    mem[7522] = 8'h00;
    mem[7523] = 8'h00;
    mem[7524] = 8'h00;
    mem[7525] = 8'h0e;
    mem[7526] = 8'h80;
    mem[7527] = 8'h07;
    mem[7528] = 8'h0e;
    mem[7529] = 8'h07;
    mem[7530] = 8'h8e;
    mem[7531] = 8'h07;
    mem[7532] = 8'h1c;
    mem[7533] = 8'hff;
    mem[7534] = 8'h0f;
    mem[7535] = 8'h1c;
    mem[7536] = 8'h70;
    mem[7537] = 8'h3c;
    mem[7538] = 8'he0;
    mem[7539] = 8'h71;
    mem[7540] = 8'hf8;
    mem[7541] = 8'h01;
    mem[7542] = 8'h38;
    mem[7543] = 8'he0;
    mem[7544] = 8'h78;
    mem[7545] = 8'hc0;
    mem[7546] = 8'h01;
    mem[7547] = 8'h00;
    mem[7548] = 8'h00;
    mem[7549] = 8'h00;
    mem[7550] = 8'h00;
    mem[7551] = 8'h00;
    mem[7552] = 8'h00;
    mem[7553] = 8'h00;
    mem[7554] = 8'h00;
    mem[7555] = 8'h00;
    mem[7556] = 8'h00;
    mem[7557] = 8'h0e;
    mem[7558] = 8'h80;
    mem[7559] = 8'h87;
    mem[7560] = 8'h0f;
    mem[7561] = 8'h0f;
    mem[7562] = 8'h0f;
    mem[7563] = 8'h0f;
    mem[7564] = 8'h9e;
    mem[7565] = 8'h07;
    mem[7566] = 8'h0e;
    mem[7567] = 8'h1c;
    mem[7568] = 8'h70;
    mem[7569] = 8'h78;
    mem[7570] = 8'hf0;
    mem[7571] = 8'h70;
    mem[7572] = 8'hf0;
    mem[7573] = 8'h01;
    mem[7574] = 8'h78;
    mem[7575] = 8'hf0;
    mem[7576] = 8'hf0;
    mem[7577] = 8'he0;
    mem[7578] = 8'h71;
    mem[7579] = 8'h00;
    mem[7580] = 8'h00;
    mem[7581] = 8'h00;
    mem[7582] = 8'h00;
    mem[7583] = 8'h00;
    mem[7584] = 8'h00;
    mem[7585] = 8'h00;
    mem[7586] = 8'h00;
    mem[7587] = 8'h00;
    mem[7588] = 8'h00;
    mem[7589] = 8'hfe;
    mem[7590] = 8'h9f;
    mem[7591] = 8'hff;
    mem[7592] = 8'h07;
    mem[7593] = 8'hff;
    mem[7594] = 8'h07;
    mem[7595] = 8'hff;
    mem[7596] = 8'h8f;
    mem[7597] = 8'h07;
    mem[7598] = 8'h1e;
    mem[7599] = 8'h1c;
    mem[7600] = 8'h70;
    mem[7601] = 8'hf0;
    mem[7602] = 8'h7f;
    mem[7603] = 8'h70;
    mem[7604] = 8'hf0;
    mem[7605] = 8'h01;
    mem[7606] = 8'hf0;
    mem[7607] = 8'h7f;
    mem[7608] = 8'hf0;
    mem[7609] = 8'hff;
    mem[7610] = 8'h70;
    mem[7611] = 8'h00;
    mem[7612] = 8'h00;
    mem[7613] = 8'h00;
    mem[7614] = 8'h00;
    mem[7615] = 8'h00;
    mem[7616] = 8'h00;
    mem[7617] = 8'h00;
    mem[7618] = 8'h00;
    mem[7619] = 8'h00;
    mem[7620] = 8'h00;
    mem[7621] = 8'hfe;
    mem[7622] = 8'h9f;
    mem[7623] = 8'hff;
    mem[7624] = 8'h03;
    mem[7625] = 8'hfe;
    mem[7626] = 8'h07;
    mem[7627] = 8'hfe;
    mem[7628] = 8'h87;
    mem[7629] = 8'h03;
    mem[7630] = 8'h1c;
    mem[7631] = 8'h1c;
    mem[7632] = 8'h70;
    mem[7633] = 8'he0;
    mem[7634] = 8'h3f;
    mem[7635] = 8'h70;
    mem[7636] = 8'he0;
    mem[7637] = 8'h01;
    mem[7638] = 8'he0;
    mem[7639] = 8'h3f;
    mem[7640] = 8'he0;
    mem[7641] = 8'h7f;
    mem[7642] = 8'h70;
    mem[7643] = 8'h00;
    mem[7644] = 8'h00;
    mem[7645] = 8'h00;
    mem[7646] = 8'h00;
    mem[7647] = 8'h00;
    mem[7648] = 8'h00;
    mem[7649] = 8'h00;
    mem[7650] = 8'h00;
    mem[7651] = 8'h00;
    mem[7652] = 8'h00;
    mem[7653] = 8'hfe;
    mem[7654] = 8'h9f;
    mem[7655] = 8'hff;
    mem[7656] = 8'h00;
    mem[7657] = 8'hf8;
    mem[7658] = 8'h01;
    mem[7659] = 8'hf8;
    mem[7660] = 8'hc3;
    mem[7661] = 8'h03;
    mem[7662] = 8'h3c;
    mem[7663] = 8'h1c;
    mem[7664] = 8'h70;
    mem[7665] = 8'hc0;
    mem[7666] = 8'h1f;
    mem[7667] = 8'h70;
    mem[7668] = 8'hc0;
    mem[7669] = 8'h01;
    mem[7670] = 8'hc0;
    mem[7671] = 8'h1f;
    mem[7672] = 8'h80;
    mem[7673] = 8'h3f;
    mem[7674] = 8'h70;
    mem[7675] = 8'h00;
    mem[7676] = 8'h00;
    mem[7677] = 8'h00;
    mem[7678] = 8'h00;
    mem[7679] = 8'h00;
    mem[7680] = 8'h00;
    mem[7681] = 8'h00;
    mem[7682] = 8'h00;
    mem[7683] = 8'h00;
    mem[7684] = 8'h00;
    mem[7685] = 8'h00;
    mem[7686] = 8'h00;
    mem[7687] = 8'h00;
    mem[7688] = 8'h00;
    mem[7689] = 8'h00;
    mem[7690] = 8'h00;
    mem[7691] = 8'h00;
    mem[7692] = 8'h00;
    mem[7693] = 8'h00;
    mem[7694] = 8'h00;
    mem[7695] = 8'h00;
    mem[7696] = 8'h00;
    mem[7697] = 8'h00;
    mem[7698] = 8'h00;
    mem[7699] = 8'h00;
    mem[7700] = 8'h00;
    mem[7701] = 8'h00;
    mem[7702] = 8'h00;
    mem[7703] = 8'h00;
    mem[7704] = 8'h00;
    mem[7705] = 8'h00;
    mem[7706] = 8'h00;
    mem[7707] = 8'h00;
    mem[7708] = 8'h00;
    mem[7709] = 8'h00;
    mem[7710] = 8'h00;
    mem[7711] = 8'h00;
    mem[7712] = 8'h00;
    mem[7713] = 8'h00;
    mem[7714] = 8'h00;
    mem[7715] = 8'h00;
    mem[7716] = 8'h00;
    mem[7717] = 8'h00;
    mem[7718] = 8'h00;
    mem[7719] = 8'h00;
    mem[7720] = 8'h00;
    mem[7721] = 8'h00;
    mem[7722] = 8'h00;
    mem[7723] = 8'h00;
    mem[7724] = 8'h00;
    mem[7725] = 8'h00;
    mem[7726] = 8'h00;
    mem[7727] = 8'h00;
    mem[7728] = 8'h00;
    mem[7729] = 8'h00;
    mem[7730] = 8'h00;
    mem[7731] = 8'h00;
    mem[7732] = 8'h00;
    mem[7733] = 8'h00;
    mem[7734] = 8'h00;
    mem[7735] = 8'h00;
    mem[7736] = 8'h00;
    mem[7737] = 8'h00;
    mem[7738] = 8'h00;
    mem[7739] = 8'h00;
    mem[7740] = 8'h00;
    mem[7741] = 8'h00;
    mem[7742] = 8'h00;
    mem[7743] = 8'h00;
    mem[7744] = 8'h00;
    mem[7745] = 8'h00;
    mem[7746] = 8'h00;
    mem[7747] = 8'h00;
    mem[7748] = 8'h00;
    mem[7749] = 8'h00;
    mem[7750] = 8'h00;
    mem[7751] = 8'h00;
    mem[7752] = 8'h00;
    mem[7753] = 8'h00;
    mem[7754] = 8'h00;
    mem[7755] = 8'h00;
    mem[7756] = 8'h00;
    mem[7757] = 8'h00;
    mem[7758] = 8'h00;
    mem[7759] = 8'h00;
    mem[7760] = 8'h00;
    mem[7761] = 8'h00;
    mem[7762] = 8'h00;
    mem[7763] = 8'h00;
    mem[7764] = 8'h00;
    mem[7765] = 8'h00;
    mem[7766] = 8'h00;
    mem[7767] = 8'h00;
    mem[7768] = 8'h00;
    mem[7769] = 8'h00;
    mem[7770] = 8'h00;
    mem[7771] = 8'h00;
    mem[7772] = 8'h00;
    mem[7773] = 8'h00;
    mem[7774] = 8'h00;
    mem[7775] = 8'h00;
    mem[7776] = 8'h00;
    mem[7777] = 8'h00;
    mem[7778] = 8'h00;
    mem[7779] = 8'h00;
    mem[7780] = 8'h00;
    mem[7781] = 8'h00;
    mem[7782] = 8'h00;
    mem[7783] = 8'h00;
    mem[7784] = 8'h00;
    mem[7785] = 8'h00;
    mem[7786] = 8'h00;
    mem[7787] = 8'h00;
    mem[7788] = 8'h00;
    mem[7789] = 8'h00;
    mem[7790] = 8'h00;
    mem[7791] = 8'h00;
    mem[7792] = 8'h00;
    mem[7793] = 8'h00;
    mem[7794] = 8'h00;
    mem[7795] = 8'h00;
    mem[7796] = 8'h00;
    mem[7797] = 8'h00;
    mem[7798] = 8'h00;
    mem[7799] = 8'h00;
    mem[7800] = 8'h00;
    mem[7801] = 8'h00;
    mem[7802] = 8'h00;
    mem[7803] = 8'h00;
    mem[7804] = 8'h00;
    mem[7805] = 8'h00;
    mem[7806] = 8'h00;
    mem[7807] = 8'h00;
    mem[7808] = 8'h00;
    mem[7809] = 8'h00;
    mem[7810] = 8'h00;
    mem[7811] = 8'h00;
    mem[7812] = 8'h00;
    mem[7813] = 8'h00;
    mem[7814] = 8'h00;
    mem[7815] = 8'h00;
    mem[7816] = 8'h00;
    mem[7817] = 8'h00;
    mem[7818] = 8'h00;
    mem[7819] = 8'h00;
    mem[7820] = 8'h00;
    mem[7821] = 8'h00;
    mem[7822] = 8'h00;
    mem[7823] = 8'h00;
    mem[7824] = 8'h00;
    mem[7825] = 8'h00;
    mem[7826] = 8'h00;
    mem[7827] = 8'h00;
    mem[7828] = 8'h00;
    mem[7829] = 8'h00;
    mem[7830] = 8'h00;
    mem[7831] = 8'h00;
    mem[7832] = 8'h00;
    mem[7833] = 8'h00;
    mem[7834] = 8'h00;
    mem[7835] = 8'h00;
    mem[7836] = 8'h00;
    mem[7837] = 8'h00;
    mem[7838] = 8'h00;
    mem[7839] = 8'h00;
    mem[7840] = 8'h00;
    mem[7841] = 8'h00;
    mem[7842] = 8'h00;
    mem[7843] = 8'h00;
    mem[7844] = 8'h00;
    mem[7845] = 8'h00;
    mem[7846] = 8'h00;
    mem[7847] = 8'h00;
    mem[7848] = 8'h00;
    mem[7849] = 8'h00;
    mem[7850] = 8'h00;
    mem[7851] = 8'h00;
    mem[7852] = 8'h00;
    mem[7853] = 8'h00;
    mem[7854] = 8'h00;
    mem[7855] = 8'h00;
    mem[7856] = 8'h00;
    mem[7857] = 8'h00;
    mem[7858] = 8'h00;
    mem[7859] = 8'h00;
    mem[7860] = 8'h00;
    mem[7861] = 8'h00;
    mem[7862] = 8'h00;
    mem[7863] = 8'h00;
    mem[7864] = 8'h00;
    mem[7865] = 8'h00;
    mem[7866] = 8'h00;
    mem[7867] = 8'h00;
    mem[7868] = 8'h00;
    mem[7869] = 8'h00;
    mem[7870] = 8'h00;
    mem[7871] = 8'h00;
    mem[7872] = 8'h00;
    mem[7873] = 8'h00;
    mem[7874] = 8'h00;
    mem[7875] = 8'h00;
    mem[7876] = 8'h00;
    mem[7877] = 8'h00;
    mem[7878] = 8'h00;
    mem[7879] = 8'h00;
    mem[7880] = 8'h00;
    mem[7881] = 8'h00;
    mem[7882] = 8'h00;
    mem[7883] = 8'h00;
    mem[7884] = 8'h00;
    mem[7885] = 8'h00;
    mem[7886] = 8'h00;
    mem[7887] = 8'h00;
    mem[7888] = 8'h00;
    mem[7889] = 8'h00;
    mem[7890] = 8'h00;
    mem[7891] = 8'h00;
    mem[7892] = 8'h00;
    mem[7893] = 8'h00;
    mem[7894] = 8'h00;
    mem[7895] = 8'h00;
    mem[7896] = 8'h00;
    mem[7897] = 8'h00;
    mem[7898] = 8'h00;
    mem[7899] = 8'h00;
    mem[7900] = 8'h00;
    mem[7901] = 8'h00;
    mem[7902] = 8'h00;
    mem[7903] = 8'h00;
    mem[7904] = 8'h00;
    mem[7905] = 8'h00;
    mem[7906] = 8'h00;
    mem[7907] = 8'h00;
    mem[7908] = 8'h00;
    mem[7909] = 8'h00;
    mem[7910] = 8'h00;
    mem[7911] = 8'h00;
    mem[7912] = 8'h00;
    mem[7913] = 8'h00;
    mem[7914] = 8'h00;
    mem[7915] = 8'h00;
    mem[7916] = 8'h00;
    mem[7917] = 8'h00;
    mem[7918] = 8'h00;
    mem[7919] = 8'h00;
    mem[7920] = 8'h00;
    mem[7921] = 8'h00;
    mem[7922] = 8'h00;
    mem[7923] = 8'h00;
    mem[7924] = 8'h00;
    mem[7925] = 8'h00;
    mem[7926] = 8'h00;
    mem[7927] = 8'h00;
    mem[7928] = 8'h00;
    mem[7929] = 8'h00;
    mem[7930] = 8'h00;
    mem[7931] = 8'h00;
    mem[7932] = 8'h00;
    mem[7933] = 8'h00;
    mem[7934] = 8'h00;
    mem[7935] = 8'h00;
    mem[7936] = 8'h00;
    mem[7937] = 8'h00;
    mem[7938] = 8'h00;
    mem[7939] = 8'h00;
    mem[7940] = 8'h00;
    mem[7941] = 8'h00;
    mem[7942] = 8'h00;
    mem[7943] = 8'h00;
    mem[7944] = 8'h00;
    mem[7945] = 8'h00;
    mem[7946] = 8'h00;
    mem[7947] = 8'h00;
    mem[7948] = 8'h00;
    mem[7949] = 8'h00;
    mem[7950] = 8'h00;
    mem[7951] = 8'h00;
    mem[7952] = 8'h00;
    mem[7953] = 8'h00;
    mem[7954] = 8'h00;
    mem[7955] = 8'h00;
    mem[7956] = 8'h00;
    mem[7957] = 8'h00;
    mem[7958] = 8'h00;
    mem[7959] = 8'h00;
    mem[7960] = 8'h00;
    mem[7961] = 8'h00;
    mem[7962] = 8'h00;
    mem[7963] = 8'h00;
    mem[7964] = 8'h00;
    mem[7965] = 8'h00;
    mem[7966] = 8'h00;
    mem[7967] = 8'h00;
    mem[7968] = 8'h00;
    mem[7969] = 8'h00;
    mem[7970] = 8'h00;
    mem[7971] = 8'h00;
    mem[7972] = 8'h00;
    mem[7973] = 8'h00;
    mem[7974] = 8'h00;
    mem[7975] = 8'h00;
    mem[7976] = 8'h00;
    mem[7977] = 8'h00;
    mem[7978] = 8'h00;
    mem[7979] = 8'h00;
    mem[7980] = 8'h00;
    mem[7981] = 8'h00;
    mem[7982] = 8'h00;
    mem[7983] = 8'h00;
    mem[7984] = 8'h00;
    mem[7985] = 8'h00;
    mem[7986] = 8'h00;
    mem[7987] = 8'h00;
    mem[7988] = 8'h00;
    mem[7989] = 8'h00;
    mem[7990] = 8'h00;
    mem[7991] = 8'h00;
    mem[7992] = 8'h00;
    mem[7993] = 8'h00;
    mem[7994] = 8'h00;
    mem[7995] = 8'h00;
    mem[7996] = 8'h00;
    mem[7997] = 8'h00;
    mem[7998] = 8'h00;
    mem[7999] = 8'h00;
    mem[8000] = 8'h00;
    mem[8001] = 8'h00;
    mem[8002] = 8'h00;
    mem[8003] = 8'h00;
    mem[8004] = 8'h00;
    mem[8005] = 8'h00;
    mem[8006] = 8'h00;
    mem[8007] = 8'h00;
    mem[8008] = 8'h00;
    mem[8009] = 8'h00;
    mem[8010] = 8'h00;
    mem[8011] = 8'h00;
    mem[8012] = 8'h00;
    mem[8013] = 8'h00;
    mem[8014] = 8'h00;
    mem[8015] = 8'h00;
    mem[8016] = 8'h00;
    mem[8017] = 8'h00;
    mem[8018] = 8'h00;
    mem[8019] = 8'h00;
    mem[8020] = 8'h00;
    mem[8021] = 8'h00;
    mem[8022] = 8'h00;
    mem[8023] = 8'h00;
    mem[8024] = 8'h00;
    mem[8025] = 8'h00;
    mem[8026] = 8'h00;
    mem[8027] = 8'h00;
    mem[8028] = 8'h00;
    mem[8029] = 8'h00;
    mem[8030] = 8'h00;
    mem[8031] = 8'h00;
    mem[8032] = 8'h00;
    mem[8033] = 8'h00;
    mem[8034] = 8'h00;
    mem[8035] = 8'h00;
    mem[8036] = 8'h00;
    mem[8037] = 8'h00;
    mem[8038] = 8'h00;
    mem[8039] = 8'h00;
    mem[8040] = 8'h00;
    mem[8041] = 8'h00;
    mem[8042] = 8'h00;
    mem[8043] = 8'h00;
    mem[8044] = 8'h00;
    mem[8045] = 8'h00;
    mem[8046] = 8'h00;
    mem[8047] = 8'h00;
    mem[8048] = 8'h00;
    mem[8049] = 8'h00;
    mem[8050] = 8'h00;
    mem[8051] = 8'h00;
    mem[8052] = 8'h00;
    mem[8053] = 8'h00;
    mem[8054] = 8'h00;
    mem[8055] = 8'h00;
    mem[8056] = 8'h00;
    mem[8057] = 8'h00;
    mem[8058] = 8'h00;
    mem[8059] = 8'h00;
    mem[8060] = 8'h00;
    mem[8061] = 8'h00;
    mem[8062] = 8'h00;
    mem[8063] = 8'h00;
    mem[8064] = 8'h00;
    mem[8065] = 8'h00;
    mem[8066] = 8'h00;
    mem[8067] = 8'h00;
    mem[8068] = 8'h00;
    mem[8069] = 8'h00;
    mem[8070] = 8'h00;
    mem[8071] = 8'h00;
    mem[8072] = 8'h00;
    mem[8073] = 8'h00;
    mem[8074] = 8'h00;
    mem[8075] = 8'h00;
    mem[8076] = 8'h00;
    mem[8077] = 8'h00;
    mem[8078] = 8'h00;
    mem[8079] = 8'h00;
    mem[8080] = 8'h00;
    mem[8081] = 8'h00;
    mem[8082] = 8'h00;
    mem[8083] = 8'h00;
    mem[8084] = 8'h00;
    mem[8085] = 8'h00;
    mem[8086] = 8'h00;
    mem[8087] = 8'h00;
    mem[8088] = 8'h00;
    mem[8089] = 8'h00;
    mem[8090] = 8'h00;
    mem[8091] = 8'h00;
    mem[8092] = 8'h00;
    mem[8093] = 8'h00;
    mem[8094] = 8'h00;
    mem[8095] = 8'h00;
    mem[8096] = 8'h00;
    mem[8097] = 8'h00;
    mem[8098] = 8'h00;
    mem[8099] = 8'h00;
    mem[8100] = 8'h00;
    mem[8101] = 8'h00;
    mem[8102] = 8'h00;
    mem[8103] = 8'h00;
    mem[8104] = 8'h00;
    mem[8105] = 8'h00;
    mem[8106] = 8'h00;
    mem[8107] = 8'h00;
    mem[8108] = 8'h00;
    mem[8109] = 8'h00;
    mem[8110] = 8'h00;
    mem[8111] = 8'h00;
    mem[8112] = 8'h00;
    mem[8113] = 8'h00;
    mem[8114] = 8'h00;
    mem[8115] = 8'h00;
    mem[8116] = 8'h00;
    mem[8117] = 8'h00;
    mem[8118] = 8'h00;
    mem[8119] = 8'h00;
    mem[8120] = 8'h00;
    mem[8121] = 8'h00;
    mem[8122] = 8'h00;
    mem[8123] = 8'h00;
    mem[8124] = 8'h00;
    mem[8125] = 8'h00;
    mem[8126] = 8'h00;
    mem[8127] = 8'h00;
    mem[8128] = 8'h00;
    mem[8129] = 8'h00;
    mem[8130] = 8'h00;
    mem[8131] = 8'h00;
    mem[8132] = 8'h00;
    mem[8133] = 8'h00;
    mem[8134] = 8'h00;
    mem[8135] = 8'h00;
    mem[8136] = 8'h00;
    mem[8137] = 8'h00;
    mem[8138] = 8'h00;
    mem[8139] = 8'h00;
    mem[8140] = 8'h00;
    mem[8141] = 8'h00;
    mem[8142] = 8'h00;
    mem[8143] = 8'h00;
    mem[8144] = 8'h00;
    mem[8145] = 8'h00;
    mem[8146] = 8'h00;
    mem[8147] = 8'h00;
    mem[8148] = 8'h00;
    mem[8149] = 8'h00;
    mem[8150] = 8'h00;
    mem[8151] = 8'h00;
    mem[8152] = 8'h00;
    mem[8153] = 8'h00;
    mem[8154] = 8'h00;
    mem[8155] = 8'h00;
    mem[8156] = 8'h00;
    mem[8157] = 8'h00;
    mem[8158] = 8'h00;
    mem[8159] = 8'h00;
    mem[8160] = 8'h00;
    mem[8161] = 8'h00;
    mem[8162] = 8'h00;
    mem[8163] = 8'h00;
    mem[8164] = 8'h00;
    mem[8165] = 8'h00;
    mem[8166] = 8'h00;
    mem[8167] = 8'h00;
    mem[8168] = 8'h00;
    mem[8169] = 8'h00;
    mem[8170] = 8'h00;
    mem[8171] = 8'h00;
    mem[8172] = 8'h00;
    mem[8173] = 8'h00;
    mem[8174] = 8'h00;
    mem[8175] = 8'h00;
    mem[8176] = 8'h00;
    mem[8177] = 8'h00;
    mem[8178] = 8'h00;
    mem[8179] = 8'h00;
    mem[8180] = 8'h00;
    mem[8181] = 8'h00;
    mem[8182] = 8'h00;
    mem[8183] = 8'h00;
    mem[8184] = 8'h00;
    mem[8185] = 8'h00;
    mem[8186] = 8'h00;
    mem[8187] = 8'h00;
    mem[8188] = 8'h00;
    mem[8189] = 8'h00;
    mem[8190] = 8'h00;
    mem[8191] = 8'h00;
  end

  wire [13:0] addr = {y[7:0], x[7:3]};
  assign pixel = mem[addr][x&7];

endmodule
